

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
BQQ8tgeoshfIj7ccAC/Rh4J85tXX6oQ0vQbmtaeTlo9mMBbO+oHsR2n3l9zvayl04A39a6l95JcW
oxkqXxvALg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
WKiRlOY4lw2QZRQyPEjgYBHF1Vjkh9uAl3uKslIKFfsM198uDcirWsFuRLqu47yWx9k/9byybclq
V/4tzvihslK8gc9ZvygVcR6dIRTZAj3JdROOVu9SueffJ6JelvF2gO7cMp61lDPW1FL5ikrO+pYZ
wensUvEo2p4nPzF2Cvw=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ylpWz/XdUZbtAmW/oqRRRgKKI7A2ZM+LZ0nNbhMN1/FKQ3mOyhbUfffJizgovZBJ92Qc4R+d6e6U
jWV9DhEXxVR37uqotk7F0AADn/iSMiNgITpgcpJQrry4XVGXU7U8wkiwv4fa6EOBd+kX1qrnULd6
HKIJOGu+iwuj2jHQhvE=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FRtTkSPlvMSYF5Q8IpWplawulFIR4PQ0aU7PUCIdf3wjAAsUUKafyrh1rhmTVaW+3nooMIT5l8AK
Ki1HVUVRNTFwoYcApRXMHs4kayCmy/jIp9PCx8ZmT9gif7ToKzhEB6MGxqcIMFBGMVgF1EC2sFJf
NjGqZwKJ49F+5NVbGt6etJx/YFXwosqbd8j95+iCA2wNMMo1kn0lk9M5wAL2v+AyX6vo4HP1WLUM
0mFS0nQsWAzyFMxm7eMd2mPJ9uQZk2SOGcVN9d1PsSiSD4PmNxEkosScepxHLbDYgYBuA9cvt9H9
n08p6Zgt6nnaBDTY6vCaDQPStkw8apPTn81gPg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
f+wUi8G3mKim71Eyhve+vM/14Ni+75ArVj1wlQq1Q1Nfl+tSD9i5FqrmGycQZNIAIg9w2XF3FJ5p
DjD/qX70w8i5nHDwjrIMxdj/CrNv/a42wBcMhDParAYGJxwrQDxKi0keAAMpdD8YS13HlSGrq1qA
zI1Ek3XwMzLxGtsm5Sr9m/DyNgLMXfl4mVH3WcpBzUN40+v/yOUHNLpkLC6P/2FsrwGvNp11l3t8
g3o95ezf5OuV41VRTQr4byMvWN1g6pNk1/EzVxSF2IB3ZVv4WC0K9FWT88Tr0upokk39pIdDBfdw
BknTcIMrJeLk03/3snAVUNRVDSycCXBI8pXODw==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ecA/NYoZ0wvyuk7d6nwrQULMS/vZZJ/1iGv3Ngw9Bc1yCpQBbqARO1NLIvGtpJOnsmmjeolioiiU
B9mksJToq1fo3rwRcigFlvjI07s7bsSvnCYbi87vzg8dq+DAfidb0wRxU0GX3hdnUIU4PB6cMkuk
028RySt7u9bGqBSXum1+I4r8HtOIUlC4u8RAvJiQ9JjYP5CmPO2/oHTeVBUGL4Ud199iQzXlms+L
BUfANMQeN2/sAxCKEuTLtdJ1l3M+rr0WOtWWQFRZDoQgZnaeVUniwCKYufnyFCadF/RtaEmaGk4I
pY/H0hXxZPr7Kge1BboMuqrVTtZT94vgvoVdLA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 867136)
`protect data_block
gu28gVZYQvux4w6FTJ7mDlqQUEqcmNTAoUu3nLny+/xyQjiFCvUW8DE3/SLYmmSNxg6GL7GDxhPy
242WaHvhRMIb5b8tOlGMAd3m7Wwho/NPKwikM6ARSR2+s7+avEhYgk1+fuLQ3yMVjgGpuI/49/4T
GEmF5jcZdy1mGUQlP5ctBizkab+nO8gaF7WX3QllMob7TnrOYkJHK3+UXe1NvihlGshR399l26zg
9IIRT9ERp1bIopnPq8GRnD6jgjKYSrEpvYIBVaECU5FNCpQcuB/CYh1oOZH4t13tqlGDQa7M6Try
qefwQ51gOmpOm2i6CEdsET5ftnDTHaTP13y5Y6e0rVOCWTT91pibTMBYgarDxQUWH5DhKnj++OvP
sNb/HIKGFyzv+cHTRp5EhdEmXIXENs2o7cHL1LldJtIh1r0VU13DiFiENjGPuGkl5geRsgCkPjSB
PegwRFolwrKY/UG2NczFcrvfyguaf3mndcpsOmKcJctK0v/b1ofJ0mK4Xd+V9vPd8LIywNI8Q/uq
4YT96+ajSwTmMpRG5ymrlsREsWydWccllBRBa2UqdQI7Ai7oKo0gE4/E/rkDQe3KP91VWzKOGr6i
26gOzFCau1LCQ0RLd4KxwlQ0CL9Z73cBmnMYjjOv44dsXg+OYIJoLUnXLcHyVaoi8SAdObUD4//y
ad5jpSgq77gunk/gCsbE3uO72YL58LKbLBbnbuKkOqfrhA6wHEwJtv+M74h9zpKFj3cap0lIia+y
3lzobeNynBTolJrPyx2bIrmp5FmnbKXRFc4BRPltZKNyGct3WXC0Bjp+YOK8hM5PgFiVY5yr0Yqb
AU5zuDNlxzj75IxHJLyj67kPBQBPNtr6oQfrfSLVX1c2+C6tRZTfv7E+lsRceb6DRqw54MWi7Khm
Nyt7tua8tfreWvIiKN/ohkuReb2/OHi8KQk3ejstFY0O32hX5KsbNI5Fb/DNHfL5Ey//DdOO1sfE
8seO1f2QFqH7lG2CRsNzCJu0ajxb7ma83s3T+JOqcH1jq1xJM0hbW4DfS1iyjJIfCVidKPCP9gDh
1WyfW1UhjCSWsWF0+AhfAP/gB6P2FzK7RC8NkIeV220daEwgwmkDRKRXeomQkH64+LPJco01YYa4
1MJ7cz1Rof23ATUmuaBsjVf36OEtlnyfFOT8M9Cv0SWUKWGjMlM8BxmmjZL4JekGG4mSyr6jHaPF
PsXPW7Wt1TYAnZ06AqkNqm+jFlPtYKLvqIY8Cax2KTIxGQ/Puj7Vqp19MxuB2ETIsDUHapjGURfu
e3i6GXCXRCkAtAgP2/VqZIHd5nOWP+LQw/7Bzr7oWNd4jwlaGlfFKU3lZT4TvJ3RdQk9KCH0/eg/
cRUfiU5cdMUB+4nLRiIHPXPRyKb/on3YxHgpjAsyBM5Jjp2Kqkdrpr79WfXlYWJ2Q3mwHaTUbKih
p2qtVejGicEqpEtn7unvlHOJUOrFcccPoHAauBNxlx9ewha4SewPWD3FW9CEr0/Lj5YhP/VV4rdb
IFwhSEf0NlSuzNVWyC0y66azcWIdEsiYsPS9yGjmMhtVgr3cX0wudLDeygSexipWqVXym6kUAdiU
ZjUEKDhzhxuZBIYLjNsh1SNynKfBPgVYp+3GSS0Wyqi79ZK8V0nLHRdtkhQOGacjr1fSoHub9sXF
gKWsjHa1wHLc35romnMeH68vY0lG/VQAKf6gs3LYLBFNyJnsgWzOF7lDjXRWja7l+aLeKWgWiA61
HSbKbTAydHwCGArgNx5xiM6rqQxILQ7C39Pi8w5h8SEzY9uSFAL8zQihWxiAP/M1hmXfyqteh3ce
52gvweu92Tv+kqT1xaVb8vLFyb+PLuLRerGwdKMresZMrfw1yBqjh/Jn7hS38VuOfOonPFNej9dJ
mYt25dDHeMUeo0B6BuS0+k/NyyFJbs3yiX4VFohkDNXnSbqWQmHxqGBy7j23FvtcZQBOWnXZ2kW0
BG27zbIUkL6hCxq16Sj5Gj+vvhR/gkeNhHrLEamDV5KZ6/rZZMo5n0i9v6CDB9KwWWSXnM8ylu2i
RQsuu2KxthqNVzS4rl7aLVU/fQjTBp/7DwWdsWsRjITa+alTtyts5eYRUg3zS+5vv6NiyOpdk0Pb
fdJO+YtE0xSAl0nTdJbKZD9FoACkwbFwUIUAOSGObiFiCKt+K/uMvtK1ergvC6qUJc1mhJwh2Vit
Xn2+zlGaaTLc9zGl+1U6TuisURjSrG6hAMrMGILFYuVI6VSl9R7cMO6D6W91dqY2oR6vWELRpzvN
l6JY9yfIrEnGcxJn0x1dmV4ZGSfhq7ggU51GLAlb9TV36yPt9j9FuIWaQHavGGl6qwNRq6Mru2SH
6RyohCcbJMTiSEWkTKm87Hr/3IhvvnpfjCtf1i3gEBR9R9YOkAA6CQgTGFlhvxqqwLd34uhG83zs
Bz2n+GdD6kPfA6edCRn1S4XY5qp68jJQkrImTi27UzKC5FlMa56+7KEVIAEasjKvajswu1LXHBR6
op8IH8iY2ib5gwUga6aX1tvkmdlobJkyK/zAex3Sz5RmMsIsKYI1/OYt0k8UDcDZrA7s0F6k/7vW
TzzLa9AwEOBuT8OluRbZi0wfGrouvrMlSuAamlXuNGJimnlm2at45nLMW/UH6XeUoh+CrZhATMc5
GPvXv2Rn+OPowEtfy3dOI0C1rGJNIwEO/MmAgIE8rQtOGLGJ/lyMID494n+TmNmdGVDODSKFGvRx
NXp35XJI/qK4SinwJ0dD+VmEK5TUfmtP/s2leC0AqXSa68klxU9ZKlcU1xn31JMoXG9A0yPKL+p8
mBj+S5IvDS4bHxCT4YH/6IiZz1kvTOlbKXzjQi3SF7zkTYbksvaJZJYQ4XjtRz64wVDza0vnrZuo
nv7o8hd4sGqE8cVMLF6isDAAt2ZhtOCLb3n88sidcCD6f54r/+RQ1axg+JslPQYtS5h6bNmgnJXQ
qUPwx10Qp2qYPLhGWhX36MYiE8vx9SJ4Ps+h8VKAzV61c25w9+MTsno3KBWeXf8HVPC6C2idvx/Q
2coO+FrDl6LGynvnzxeUEZfedZUFD8qDfpgOvq4dcatHI/s1mAm2e5Q8/RdP2nVHwANRIYkk+gjD
FOwNI516yqCBLuuKPSjWAulGnGGFTzdujvwLpznquPoRZSSkA8qjlpPiUWgPoL+lsLjsHewWusAP
xdlhEZZC914NoT4DJrzrXGucIbg6hKS1adMZzdQQKsaiadPFzEXA27lo1H0PnPFcUCTocc+yHc9C
BUniMxAbNrp4IKdaGBih/iMquRWE11nXg056SFzvtnW2TxhRGLakbElkXeDVCcQCSEvXhiJSjiY7
2LZh8T4lyMBTF0xulcdLKLp9MDUuZNCZ3hd29pPxajECsaZ6JfsO/kiXOua0Sl1dcCS5F7pDE6Wm
swfAyCyfX+r4bBKOA9SrSkaWhcqNFqzjdXWygETmI5NiC/Up1qorRpPMIfIw9R7z8RENHseLT/Vd
rxonbjrvXjdRzSJQV0IxPA8K5cNM7Yu4p9rxssp3qQI3rLK7meXHz4QBmY0wE5bMI/nio+vs+qdO
AiWlIvM71b31I4evbnTSr8kkFQo3hsmE0CAN5x55dM5v4EZzxzlEaJnIWrS6FH72BHBP8zSqHHMA
fUuzMOqeSJwwlrjviHpMVBp5T3IwYcxTfvSZpgQCYzX8yFa4GqG6v3tWdQBLSiKQdTYcM7eAuEKh
CPvU8KNYIJIgAWPNEAs4UDwjJnW0zZuRbQnMt1SXjrHM3G+LLUmqzxDFQytdV3kLbQvI68qBUylw
wOlpfMDLXy5CRDUPybFSWSiCTfiTRRBRG1u7tYXCYblx27pCdQwcmpLrTS9LagunKG+mhFtk2D/O
PEdHOeebJaWj4ORvRbFnAndMaM2yuzx9GfjVRVK8ae84rlB8XpdaFW3gT6tclbvwjOIIjKLthf/g
khpvnYFzNkIBkR9xTArZ6cdQAhbY19Omf6lqStb+099qv51KTIcKb3ccM1NB5X0LVXdebjYc8yRi
mIb+5rcwf6y5IBgKBqtqCnAHHNikPNKdDBJggb5sCvAadoUbJkSQt/M2PfzZ/BmiX585WuIrlByQ
wninZWud1WwRZq8z0r6VhJD2N4JIszKKIWiAVqHb8h22x6rIxJmOpSyyY+WFhtbdNhkLM8FtUUPC
DtCG/p7WJBDo7g50r/lCi09ToW2bht4N63MojXjAsU5VhfAk3DeJH9p+SF1XEMpldO7WKxQSQfhS
3dKDw8aeapg1pvh6QyVIRbo97dIqdEkn61klTbukyESfokdPjzW9rdzjKsRwkPF6NyrPxVBnCWZ2
CXPZfqnLpsDqozb91aF4uIKJ477W9fIVVdkNu4ikmSRHtdmJFlUm1peQxWqxV6VEkCCvow/beZzL
MHllAZdWJNWb2XhSKbxdY8FncPuJPl8EnIk2HAmZ9pLtqjWCJlNrU8P7PHrCayIrRg3j1EN9WI0c
tUB5pAIsIcOgQSnJ9jgK7qTlONrDIkzE1VlIBfpotH2SN9eZduH5MmhXFKslqm2qsV4Et2RuSN/O
C9rvm0XPlMRcoFFPcdKrxG2sVNk06+faKYfHPptasBS0NxDv9mXXPh5hRL+GD/oVA1tsBFi4QjdQ
iY9HkcaALjNGR3/fKFMOo4rRHWAerHkzZ8s5IOanJLJ0kdkCVn9tZgW4Bu43ug0lblYNHxZaShuz
2GqbgqltAPZNaaymEPlldCctfE4UcC/ISjlKMqBpXZ0bnHJhqLY/g2DmMjMZCsCUSa5TFNJlU5hi
uczEea0ue7ChoEBxYouDcsYr9bCpWq5KNQYp5iMYjBL/z6fdQq+xx+zp46JHU5uHdVA1EltErZSt
Y2zasFlE6Mb16vMJvzFUDNX8DNMHS72Dfii7zZuwzH4FMXPko45MjaqLzVAlma9lLZQeEUr3GEHd
wso0zhs2dU4B5GQd9onHG1q4bLVMYmIbMERhYTBdczZbaAg0COuIOmrLCdg83IfSCrlmQWeyzgRl
pB4Mc4/yZ5jNiuDZJepNvsfWeP8t2lBTUfmP8gJyvvlOOtjJ9lNnyUe+eu/nRLOCws06j18CXuvP
cNZjBTVbg1l/qc9eDsPLZqui0sbieUDwdGCa5VvlEdLk5Z8ITEs+IyQQS+KPpbLNe3WehXBrwsHX
QCg0QjfgfsS8lZOzNStkmGhn87jAJQruQfhg715RGRAOpFq/RmyGcwBXds8t7Uw0N7oCxGwTZYMx
6wBOpqxUmbYlbUIDtgiCq/yeuy4SSy5Rhy3cgJ8PSHJmwWNf92oNRz5sR7byq4zuxc7RdNWAtchI
oasCXpD3EDW+WruMju/4SLWC++VA0aCQDIahos9pRmbnvArKsH1HD+m4nCZXqLF9YnCM8Nr4IANE
hhym5j1dspvzeEdX6zGNB+/EIH/MMUcT7oLCZCq5qS5pUIaFFB170XhLvWN5T9Dq5vWvH8Mk16pS
A+3EtrxkeBWpvE2EiLPrQLAtIo0KyAcKlKoQJOU6Vq9rs1AGkqqwATBl/Jskf9+vAvJkIfl96KXH
XUUFIvkCf63uPIR2lxXh8J9zxADd9xcFm4WajUHo0DZUj+ime7BxOLZrX/J74kGbcHEMCOLECJZj
oJpHfJdXyTvdSyeeVNyiEMjJQHEEQ8UKPE6nuHBG1tmf23+VCskB5xnJVMF53yVNEz+bMF09Xd+I
Dt201xjUWOG80FyqAkVQ1y4rvCoEVsinUWlFHXq3bMeiT9qcF7LH2TGu89s54lQgh2PdxClarr8P
kq2ZxBYF66j9x7B7H7DfriqyXsF15Wjk9j8btKboOXffUAZ98soy6cDtnx5BEt72Pe5dL+6nBmoM
chPmpVwi/9FEeinKzxa+M4YGlmJlhjxvWU8DftYzp0wXb5uhvG4B6DwwJVaep/rXqu5tmlqklb4d
WOiS9XlOl2hJsSJ5Q0DbQXZIYYDIbiLuxWLj9V76wCN7SSIBYr9OxqRRdgYElRDhCiimquhoetfk
eJPWkCkYLDRbxk89OR0WrQUMHbjhaSK4w/TBrkSgEDMXzOGCQ763nN1o25r08HXpyaBHfoSclzXR
cP4rA5SOC4kdutYEH5yIXtZhGyYV+ZCQzWV8KW3g8hBHmCzu6XQkwyAvpkOpCso9oluCDHTxIbyg
dnz1rjhT2dn1RZGlA3eQxxmCWxNZWp6NpOIU+HsWnnnBs9cd+3Wj6PuMceu1NoqS3BrCU1FqDyXo
fQHQ8zc41XGtLo4EG5jgXdm0iaHeIT+D0o8hIWZ7keAwPEKehE/6wFOFXkFAx2prOf+uMm0VzbQW
uvCq6/Mu5/ioboZDI/bD5w6V9FbJp4hqSHKn/PJ7vlSAaDDzQ2XTvJfOtLXa5Jr82vp+Nu35BuSY
/NIel91YZH8Fep5KgQKtXCXVUHltP31bAzmdkxzGsFvrKGcW/ZoDTQllrDD83p/bNFEnYPSehgDH
Kk6HnDhRgukLQqzSBFMj8iH3snimxd35zbJP9YTBin92hQsUsRDuQU9gEL/jB5PTZovig92x6Nc9
jsBaS/oa0SpYi5qYL4q5WfJkKGHwkXtSB869Re42wUhindmXhCZtT5bsVwIHB3sQldUthNJb7Lje
ONMq9ARz+HEXXbY7Mxl9QxvE0mBz61TrxevfAw6hkfm/28D5pi50a4YPlTI4nMktppTZ3TcryS46
2wKaxPDvXy7KBuCO8jv4XkQf9SGmOYOWS0rsOVfr0efRaXAG2IOM3iqOGgoroIYHtIB9kr8eZoTV
6fk+HSIiZtXzG4u7mN26Mbq3S0EZWFIHC8zb/hRRRnTfdguaCJd1zCddH9e3jxvg7im0HmFaRqvE
vX7BnxCwbZ/ap9BtCXiTIEzBU4fR8Jtd9IsFxLYT4DLUb/7QA/8/oTljHFTaUiNaxWiMKr/nSoCV
BQSPgobFWNQ3v2pc9PmDR0+SvyIu05BQkuJCcWfPtwh++MqiBKK9npQuAGbe2ekhEI5VGRui1n+K
9OTb6iMRsbm3toZu2py8HxaXcOD19D6kccTXhaZPWF1ZjVyunyjiwj+45F5Q6LTg0RCTbZdm227V
rMcJTrHfNAFKShFlmZ4ciWpA/G15HSKRLc8VC4yDL49VWPuqgMiB2k4CP9/YBL2/JNstSH3Eqvxs
7tBOC98/7BMjz9NdmPeMXvUW7o3rLuPz6WeBTthZ+q3a1OT3H2+0dwNzbaua+Kf6vSWSm2XXbD0V
LW4J2gGmEBx80ikcXlFlhXChnEPX3AqocFAlKtqM2rVNwf4uaK2/1j7I9ez5zGZw4AT+ob1o3F6m
HgcNjQHEwKeiuioSYxr0YlfEuvchH/JuuPMnFY8XP/j/Qjz63ayk7UyYQDuxDnOu4rloW0EIv1tL
D/125+hwnHWsE2dh+Qvby4n4nzvo0diz72lSQ8IO5s9i8/HjVmfc49AyVHz/kPTxGxmAy9uZFRI8
1YySaPWGEUT0w0Vr4cradJuMhyG91s+3hLzU1YOTVhE/JM4c4oElNYyhp1ISqdM6K/UaWJQOjvKI
xQQdeDc4xhPGpd9WM17uhvEybNS0UMlY9lf5nBtUidG3BdT9nj55fJXsWkxFxivNEpsy86Uiro+t
wQYXYl2kw97ZbDRD9PvKK8Rk3qRmP2NYuRcKE9a/wN4M6UrLo1okl071jI3AWMAgk6ommHgfeeyM
ixZY2xrzB/0VdB+H/gfWQJ7sEoqi/M2MsT/qyjt/8Oui7r+KhRaSCMAwnEPV8AyYT1EBuMu2AWQk
grmix2dB2bNsIzZQdexpuXnFdesf6krzaaA6kgrFYp8N+bW2PCaEDizQRLe+kTx5FpWy+XAdLYfz
RQnmD3XxiKy6dEdET0f42e7C2ACpaRcax/wPf7iu8ibiTLA95jqErNZaK/aD2AmR0zlWH+Ax9x2X
eFYrrNFRDCXSMEasrOcYrAw64iV3UMkiQDYOpuDImsZbex76KrugjkOSlAK1C8qITMX2ZeF2iQGV
H8poLvjE8/qmmqFeE7r8MU0Xh4JSFM5CQkaWQbY9tO8ccZWTfvUhjOrRM4hngXtK2hKFlWq5L2ej
euIoptK6q+9ovdp2xk79vSotYjAmhhi/BvNd2Fnq6USgQZ0Mq+6jncXcj8bw01ddeeX1oGMpwF+H
/whcI4p16YLSLch9pJUPXZ7Tb7vneA2tgAD1j7OsLwD3I9Li4OnWZ4jDOC3QOQ0ZfIoxfRk+34W7
4yajqXvK4ZPObK/DRe+GVH82S8vIpPXj+DlK9E6bdKbp8UdOo/Zg1qHZQlV7wqqQp+rStMvrAFmr
LDIyip6dZIsRHMii+UkPx9H6IC/SGn1w+/mW2yyYE+b5fj4a160AQ2gbsKZAZIQk+yJ/FqhApkHz
slXn672tZGL/yywSlJs0+n6aZofYd85EBqW50XT+sLEDO1aWeKR/FyOLS8bk2uT6naoSs1cIutSH
Ky05t9GN/mC1EDaF0t8mqzgMO8gbu/7SWNhpF1qvjv+7azSAgcrvEHy1KOm2WY1mwvT2oGm3OnkW
W2xqgsQNlg2bGJ6su2pwpxEkKyMSweMyqSsJ18Gdvbo/vLNBJVRWbQky04dgaebLIfKpkin+1owA
0WObtfAWuc2xb43Ax4OX4vzQTNyJZZkjuifCUhTsU3owv+HNzdPSnpYUa125j0newU8EvzUVi9aS
ztQq9JTact6qK1sKOiSql92175NJVwdnZsdBX8Mt30/Z6eM1eceozQ46+cRp03rI7bxem1oKHXHm
jU51LCpDK7WWEUq8eDtFDr3hvJzfNBur52YByWBstSOOD5kfFcPdoZCuDbU2KRCPi+nk2l4GoP45
61J7pE7vv3YAKi2JzGL0yTx3qh8S/P1BJyI4ExQKR3Gn/h8csvaAG2R0S/ASD1nm4HXCoqm4oEAY
J4GYwes36j+GEN5NI4RmvAHIKkSx5pSYMYnydOExTDeuSIyOYO+RMJaaW1Xrmd3H/VySNpxdCWYT
yUSyAzXXiKCdH19L1MiPBr5v1G/sZaGj1Yof3TxwgGqXJ7XeeOoivH308Ebauw3lY5wmMHWRL5N1
GII31FqXvj3auUsSm3yNXF7LAjFCF+QhW8cVF9nfaXbOAHtmVa/8R/eeP7qqxT7KQntJTY5YRL9N
r02x/pTk+xY4dN963Jm638vj/Fi5GJJkQgXd1fMAV1MHPK9DPPWtwKe4dKvGgkReeknozOO9y5Zy
D4Lrlv5vdDm8/zJvNS9VKsvvk8cz34/73AwhMr/AbOjfa+vvIteon6nmPOOePn+mTrHfkVzcud/o
05ofCd5f/3iBGALvwBlI8lUsJVcuVQKVaQtxHfvTGAm/bvjwmQZdiMHN7o6/ROJJkd+RfKJIVNvS
EKbWjGc6MA5cemaMIe9NpU5BKfbz7LUMjxL3Ly0wX2GqBWSoXOd+thLfEntXK7dwHpPB6NuMWOdh
58tj70QUiW3TgeuP8EGaQHtKcgbVPUJJXkPhazklnu6kDwlUVLdIkkhpohC+9Qu2FNRmesJvo2R0
36t2tt9yJA1ahAB2Y58nf237GpRIZmsRgPZjgEVar5c2HWITSu74Zb0h5irx+OuEJ64/8kFX9uAZ
VETDTLLKk6FFErnpwbC9KPlsuFX9d2lz9cQlSZ/irvE8wzRhG2gouKkK3ZXwdox04xGKTpP5qirO
iJSASO2b+8PLU9+E6qBSLod1bS3ZG6L04/b6UDuN5Y14TIUmwZG5D/YUJEyqW7pAcm9e6nBu65RU
huIKbyIrbbTuo901pGaERBJpm3sZI7zFy5vpQPOyOsFNMOCyIqjp5NaGxI7FPKmaSoTwUiq6v/SG
6ZxGHd86x9J/LKc9IKs8OLbw7nxE3K7xc9yuynpPZeHGBksaON7JAcLabmZskG6XeDk4RMtTZbRj
aZjUEL2njjaz9iyBPQcAEWfB43gqdSXLIoaiL4HPUCO7iotoG4SNAIwXAZh55zqGcTgJqWlEmkDR
uOQDAKbJar8n8rMnWC54G5f3Vo0We9R4iMlm/EqG/lj7gkQ+1Dx7dny17tSD1eTfa3H3+PJralWR
5+TK6HM/ibEgDcZwQv++O6XjwQk1dWILqGhEoFr1DnFQtJd+Pz5tlVI3Z5f7xRcCKCbG63LRbXIt
fO6Nja6553h2a3Dri5/yKirho60dNk8LopD3O08tydVrqtZEUmoAocp9p2lwyhr+sRXv1sK1Psxu
MFjCrfzj/vSRoZaFaY5Oc4UvKh6cNWdJTKhTuE2Y0Ne+dxU88CkKmgfyq+wq9PulSo1w1HJEXbD1
PHjlhiihWIgik2HJxsErVFxVSMdDJqrlw4ynKAnAfV0Xd+bsfhd6VMkEdNNQa/RnZ0eJMqAteUOX
dC/sBWt+gDLxw+pYo2w/CuxUD1JBFYSx7KDl7kKJKNtbP/uj6Ru2PmcXRBNkEp8gIxgFam0v5Agy
3zZSe7kEDWFaV7yWz5Lu5sHW8+cvtxhpgyBk7MOZ6HPFSV5TM1QkvQCqpZd7y7FbViiTQJ4z+CcP
CZctDjYef2pLPO363JaOdk5r1+zniiDtz6gDakGoojtpIoyaVk60/1Pr3Gb1hqRVDxQHLixGIUrK
bB5PWxtfTxGWiQpTVzNW6MpVRufzCEsGlaYcowMuz6u4hh2NKZHeFeP39ld3EQcxZ2vjcZv12YBG
ljKiXRlezl0MmcVN/dz0OrJp/TfoTML6iMqcLtoK4vazoH7y1liNyazIhj+wUG+jkV8rSvw95385
CF6SeHxv3pbx46mU05pRRR+UDXm7+bSbxc4Xk6KpW4swSmEu9Y4ueeMEVznlR83E2hSd56jpkK34
w+IT1B82+F/OU0J8MCWAh1F2w4P/h8z0iyuVU/XpBfyEOyetd+UKR97uS3b7x++QQfyc8N6q9ntV
RKSku2+6I4ROCSRaQ3zg4s2oQZt1mONeaHDXbltiOTJJKL2DC1Fl/Qya42qWNVYBy0Jxsgpbgv1C
UPY7LOEzZNW37bodS5+XBYZxJBWvLjRCWqg6R6wD4+XpY9eRygR3YUp0jDMhutmAwaD4e8kaWxCj
nhBpaevx42FhHeDS+15ygIctKtAMU2o5J6WsZgYw5hEnVeqnIE56E40qWw5tSQrqaUonNgSodn+V
PV8nAzK6YE8oFqWl1cteB4hRVWQD/oNMld+Q2i5/bygJ9HY1f28KV3sqdYa8K4uL9qFEhBENOccd
v1jPypZEgT6wvHqvqgkcUZFGbgroy5+Q0fxfTKhmHuC/7LjzS0ja3EsWjGYGWcXNaFHg0hD2C/BZ
f9vPCfn3ZVp1x/u296fh76uvXdmWNqbJsLp5kThTftxPZRSGI01rRFlg6uoLLvq1IIgcXMmDtSq6
Kldl8upM7+h+jQKC0m1Sl/spFbhDb3jlvOQW5VixM9nomPfaqyhWxI07uCjNZ6V6frLcd6c/ZhQb
TuAt4KK0rtpWv508xYTq0u5C3fDws7CiTSoWXXAl7P748q66JcvP0ZolEsgx77QIJkXHAFZYBxNX
iYuwaQH+N+3jPX3suyM4P+aoy7F0WP6Xyvxi0ZuChLETstTj9pMISYvE48lhtQIosvwkJEJgRrXJ
FoDmASoZcCxcNhei2iJWZ72i30zTCgQBZbqZ/toVjUUBsum3qH5JOC/ir8+N2IppeY8uBM56WO04
2ujQKNh3VzOY8e7MwBizKhLxGGe855vzG3x7Ia+QtkYgGCYtnfrifBg4tXXYWAEG451mnghRwhJ8
C5N4x8+8D3Ko0jgMktuuumy28PjXHJsMidSXLAJbDpttbKQtP2J6pDMv/TAaEmieI3tqlpJXZlAZ
xp1imsexJUqjzC2u4ot+474PXvh/UVvMvZaMFWMITIdiKctE39UOTqYhF1XBmuF/1H4Bk5hGNIYa
4Mu3113aYWZcMyDFiowMo88BTJL/Yv0p79JMYq0KfRo9wfzJ3NSJa3/qkeV9Xl3uekEDI+xQR8eP
48hA9pCuVYvg/BkPawoGKiTe/wC0Rn36S4eVkbiIkolWtbGN1XrEwHBuT0LRK89kP6lATv2wpO0F
jEZ0syLM7wcgjqek7LZnXrPG+q8eNmc/lzWBxxjTfbA3SN34wnRq6PlPZvFuxpHrVwys9Mxs5fsq
MRAySNe8keo4iG0Mo9dCHE6E3TYwUjqu7VUxLczIvJijVpbFz+QJxH8goypGtZnKG8u2ynJ0QGF4
+FxfCqEEwXFmCCz4yQsp0txvukjijfjLil2ScysiemBB8z5aMxOGKIxi5b1+5eCyN61vPhaZPZ9y
GBIA7uGSfc/NiN17xH8VRjvlzNtRr3QQEGB/s7cmqxWlepPNMrAGs4wf6YWd7a/C1c+bsDbXTYOb
9DzcVbdBh2VNvbxgkOcwEak8nv/zuafodAW7SmOHlpRiO9CAzNEyBI6K5brq9UFR/SjW4l5Aqd0+
vejdaHXQZyP5zP6A0O5+s1FVDoY1JoLVnybbe+87omdBM7APlk6Rts3zM1CsrFUO//gFw5SsKkEK
yKQM5853JxzYFvRgVA1JDguMlLrnBcFv1fnTHDfET3UFy5n3adjgzkoAcBLzc9xL/28Bb3NjPojr
6tyzjsX8UgKtDWC9APgcrFhazU3EEkxkdF/Vp6cnstt1Ab1JTteJKZ5r53WwrRp3GBlYN8a1N/SL
GemmIZhtEALmxSMC11d2KMaw1x3FTS8srQnEI4XgQZ9cN9GdlxZSdoYRPlrjN7HmSmcBbOprS+wf
Sg9wRjnNJ2/DgcsBfLGaKI/L8s6ZSTMzF138amP6R6YJzatfwuM9+/Rj6Lqzf1DVh61tvFnQbrhG
sz1Z8hUqIKVoEioFWLz19ibEU97IpM4Ux2j/Wfs5noiKef8t4rE6of/YWSwTzcX8ZvLfWEAqm0C+
kJ6rIJMSEDATlmqrTeoi7Tb8o9X/NfUbOVVD2amI2w9ToJJYePDe3umVzvv+sDrS51HSTcQ6ikiA
ThWmWad6gc9XBpit7E2ZUXNSZylhB0vw3O63ZlJfkau2JtkXygiqYu8yEvB9Yf43Qy2xRfTMQRyJ
TL7sMVZyKFkUMLEPSJlzi9n9hpORq5zlq22kdHucwXqlhqCryNvfjH+3N3F0pZdaaHMrsHi1xP2R
S2cV3w48GIT5rhlsbeQgZoG5OS7zMOXELl2gIqU6wWVNZGXU74/dkfu14p87HVJi8iUqdOHRs6sX
TBjjIhYndq8vOq+W7gcllvPG6D537dIb3ZchXKgzmtmooNeo9MzeJOFXnYKvLKErEimYuoOR1+MN
rglP7N2eUJV8Me5w4F6mpaxQ2qGjIGGTxy/JRJjMCNsijbHQfDeyLpXPFBqjgNhgmdqPpRxh6Qm3
XfGGIV1OLQyljZYjzeaV0HL5gtYFXpWF+jf1VxpmWkVe6YOBfe5Uch/i66o4nw3xQMpWTl9DmJOr
qK3JKhf2uusTzlmQYBB0+mV3BnYodV9oq/t03hwa1AW4v4RkbvQV5Ak9IK9Pwf+SHyXNneuR7haW
tXGDkLhkfmcrqowG46jFFN0ZWmcWCPGLHyy+VC3/ODOpaV0tCgOD03CAczVTmKhz6AK6IV9ZEZzw
gv/K9bzL8nx6IcG+vOUHSbFZ2xUgt/AXi4BjF+9mNDbM+1w0z3FNwGBdSSHP3tuf7wmbbinyUdCf
iA7Vn3toIwNTwdFwolBTJMVRRIrHNltE0IR9hXSXOriMbKyUdNpRRs9rgYgccYgeuGBNRUlJVnT/
BPlw1z8w3vaNCs1iAadSxZg+xGUw8GL5fOWbnAmbzIF+GY3lGqcxqIZMLO/itkbPup+1vPOUm1TK
x5v4w+fZpM3J0uv+F90BNCkRrp4eVdZ7RXAkIYgkfLH/TJ6QX9NhgY7NeT6ZZJNp4u7Yic1Z7mrl
f/twX2PrM8o6NMfDSrSrGOf8rXDXKD83nrEU4LsPExPw/v3OJaYPqLPgw6FUzrnN0o58XTWX76qN
U+b6kSsuByMwqIbtJ/5dbY0YyVQPcgH3DyY6WM307BzR/YDV4uN1zWGyJW+/qrVTfujkV7K5uhpx
67UjcQmz8vEQPTEVVMz0FF2upqws2D7akWpyT+hhYloNpef0tAmm09HPOKk49dl2wL5RVx42uh3X
7OL2USnd2cusNXenQFJXoeFgikvFvkDu2WHlLhvETJ4yb8/jY6XxByHY2Yq2AC0t9EJKMS9Rzpfr
jtIglRTWXbJLBHODE2uGvPK/ZCrmNzBrvyLo/M9u9hO70uPeug2eSAQHnWyjVefkzFf6nZXxmOTi
8zo8pA9OAhZoMSX4PMm6FRpsgYccS/yMxbOC54MMiE3LXnAq3b8VYZjoGC6ANqkFArxV3djoDtOY
AsbhdRLakQh09Gr/Z6Z0YPofsbYC35ZJXM58ZPk7j+MR/j2/YHrfcyixcKhqMLnMShFBa+JwJbN0
jxKWpCixlUOfynEPzzxSmUrSjkXXLv3a0Vi7vy41mQjuakaHgwQMyLRYA/ZfAY8h/rZIF4rrNSHY
UXusnuo91A4B3hbFMOAnknmf8Zt59qGgCAUg2rS3TKRlwxsYXGczyjBOQSZCLirqkFTlkJUOgSaG
Mrc8n9cV8EgIs9D27GVAzwrDz6c3SG+W1j4xXURPz1lWSPUkvcUiPhF1FfASLFzfIrvfq8mnGQjJ
40gQDRt/ddt+bpHUSrEoFOI2KknvUcaDAlplXlnvj0LDOEj6mLyrCc3wcRpggnMOeODf0ddBI2FK
ftBWDv72LNdhTo1R14KH0ZLRsk4gfF+5MnomuVTxwHvvJt7zYbwYOiQ9hoUg/c1nB0j2o/Jl18U1
bEQkBVcFFj0UqMT1oURPXUWmb/sljqa/v9Qds4YRE5zxPA2prf06hC7wTS4ZqU+9U4SrVQfascVv
sbxCsCbxe5FRA3UvwlZF3T5WJg1KrWJ0fM2Y7x1M4nVV8jnQ3wP0xlaU0BTYfdZeHlW4f1E0Rtmh
/LLHUBcjTKyWGKYqGQu9hyl0DR5lltcdeSNjQ+GMtxYS2rcX8+NxBTVbr44CYksjNxwD9QIexYvN
3qrAOBsDzcozi7yWTOz+L2+LKs5TAjWIbO2TDB5UkBlYo6Ywc+CH4cAfnwKBUW4MG6EYhW7pia3W
xV1wBp+pS+bjEqpODqv4+EHQa2/QBwMZx+5TvLXCTJWKBjZrjwFfR7VxNpi2C9ENIMiptwuKhO+G
PxZICmpZIEzpLq7NMvFPt4GhzM8/aH+DBYAJolkmPOeSG0S5/SiuYJDiUedOZvKsebQJ3bGA44uw
ci9HwnXIEfNTe8oZyZOjheDzSMsxwxrfrn9ES4jVBlhw0pJbj6Bvuphgb1FR9v2mhMWC0lFPUIVN
nwbFhLN2l/Lly7iiY+RsnAO8DMxRQI0x55HXWkoaZdBU+IJoMMUYvthfEI1dc9IosE9SYqwdXyeK
SXHnNAr0++yR30clf6CpI7hPgPBJeDzeb+2By4yjmVq3uXO2w8YOXlVIC+GDYL9JwUb71ieOsye7
gJBal9kLgODqb15ANTJRppDRHHWjJTBucoRpnfK4s5e4tNlTQOpFJk+jncReOiNfBpTpe2Tr7vDm
ifdfd00J44tWiOunlIO9R4ErNCLzm8uosxnAzv8hUyVKryT3CrX76J+7v32iiawXZqfLUugf/9kQ
Xpnvs1hDAIiJvTB0liWQmxjhyNvwp6jQ1BbytN4PeFkMUXdDs9HdD+HWR+IZ9nYBsXJIw+PSG7ZG
X0rLrkel0+5fl/DNIiLEwevbMN+9FWC4sYrdB6Q44UC4rWJxRAC15DTrP+L5vMqqZuZ58JrMwWk3
UP9BI5BvbtnVs3e0I/voobRxzSd9nLKC4Yx8AFkfZiSxGcCYm4Yuz1nl6ADryBZ7XDu0kmdJxZ8i
hCQdxUZQgXZp+pD0Yg43fXobmEhb+2gkon2OVzFAuKmabGlGBJi/wjQDO/ic7kWZsBd5rPP4sl7N
HZ2+0lqRQEGPnHCjMTx0Y9uGJ9vVwDoOa5UmbqrqfwHESqxs+kJOyArK3PvrOzRl417zpfo+IPV5
TlK1B+FJuGUhd+7iVfSZvUrqwaPnjLiCD0SGtumJn0HmJVeu8QGlXOBFFZFt7NsicRpou/p7TYrR
l3fiuYC9z1UsrJk2zq0qi2+QVj8kJ7juJ+ANOSJJIrNEnAHQLsT9kZbuIzrX1OP1Dt+9u0xnkr7u
775MfFwCgq6peLKgaD2kvHTxjlSsXpCiaUYc5zNkFBaOL0PA0F9H+E6o/DsJoL4CkGcQ3/407IVE
MS8YqlkDo+SK16WTaiZFimGvqgAsGXg1psXDfVlNR8JwZb7+jzKG7LEPJ9QLh5D/jsO8SoqGK9np
1AcXS2tipeMLaZ2Gp6dTjXXPZjcdGW5CsjF2ae1yQRCVIWK5BTPbzflls+uaHJDTnzXYLjZDIAFX
ygl7491CBpPpkZrudPBHKX0dqZMqjmc1/yQGQX/QG5QkOccvZ6dfqhoRnbouboONX1PBlhUVLsDa
PU4kSVXba3pfXet22+h0BjEzkYRnEAHd77K00qUyra0RbkMQjpamO5kxB3eahIVY1X4MCjgVCW2X
pgTe9zyZVaZe6TrBdhDH1NcYHoWygCFAipJSgdP/fVnsNEekAH+E6GGOsh1M9+r5qvw51rr+gJy6
ayNtRatpBU7k8A6zq3OMoZKztRj31tr32X1DWRoMfEDdFLS/oiomWE/EBAe89oRP9IX8szlcHyNQ
dnFSC+1ypXReX5LKRaojWIShNs0Ux49xmlLLGS4SDoTMdlTTbQVT5ZsKQ16C+lrh86MPZ17rvE0C
EBLMQShgrqUghF3XyQ7mj4fQwgMXLqPeViSrA286F/U/EBMmWrSx+Fsx+lpUhBMMpfaHj1ZhnYmR
+3a8uuLAp5J90Ui+14vw9D+afpkZeV7cE3SQXiDhwMi814PWUE7RRzr/IOqAgzHRqS4UnF6Zo/1s
aPsOJ6i+9L3fx6aq5QyNJ5MWkV+Hlwfb4jK32AcEQiukr8g63vjyK2acfzrKRJLKNpnRVdgXqn2V
ad9Nn4fsZpMuz1uSLkye2UomyHhe57NsVp2C4d/F1eGo2KLYHOYcD+jhJZ5K5GghjKVAMUdt69Px
sJYaAiQ65J5uqaF9/JAykkNAWLK2YqMcMVIpfmL9Gt5sK5/hPjelXNhucX3m9kFFsQphpYzVQnhk
6rLL9kCKnUQWmwrccI4LzF6gP7ycAidx7F5kkF2yK6pmS4k2vl8mDsaaKKyd/BKED9C4r79uHjeN
bU//Dm7z2USWvijBry5Tg5AvB/OmqQfwrzIfxsygF6zDF0E2693wwIX7/sBgu+0kxqdCev2BCyL9
eq6XNS5Lk7m65bhAszaV2s6RV5FoS8N4Zh1j5Us027RzFghTamDA70cIq3shJFrdBaNRlDdpSvUi
hZCNqGJXQoiOrUWadoDfHGrf8iV4dUzd0kCfgDDEH+y7mcd6Rw6MucjS/MbOQO6DfMe75JMX1UVe
maVO514h8P9YgI0HaH5m8YFNzaHvlP6yGfntfjxmH3/4OjKDZZPP8c6Ux2l0rbFnV716QZZNAKiM
FLQ9ICuQjeLudoDnPJbtGTLYKxIoRclMdEG6QxoRaF9JH+BpP40M0X/+q8/SMS4RECxTL4CJDNiw
7jTClrzXVNekARuwf76an2nWRblE1QDz11XeG4kEJOFWazOq8WK0Py7WqHmS8m9XliIGoG1iDbl5
1ArXND8vYqGJPlNpSmEdTaDi86zEsoRIIgz+m53Wysa9i2UsEGwgZuGdvcoeAVKufyhn28uMn//T
drlaoOPuWTpLxVbOPpYkPgOz/GHhYkwVMS+UYhKLxYgpIeOuaNlhFp4jAuxi2OvfemhghmfmNw0z
1lHQ6fSQBbr43Hr7126WaSy8Q6byp5VxHFHv3v4XUfQUiiD1titWcupz1wh4/v2guOp+5tT1kDZN
QqiQTkVzfLsMOTvTHwPU5EctJHDqal3oPimZ/iGErupVKHOjmd6E3ZhOQdjQJHTOTQfMM7R10Df6
VneVzPPb720GG1uDCCA4HInteoPRYbp7fjQxEc/93HZROB4Blt6iEhWriajGVEjAoQ+GguzDNzWu
OWs6hH8SDe1B1C38Xgcd0TjzTEpwHchnsP43n/3MW38d24P+ickvN+iLG5aS4sFW5SEdPoLKlxB+
EOqHrLMQm0KDqjM/oqua1N+hmpkRd44CCEZl/nmsiVLyDGIJMTOwUIQqGzDjK0ITaiOVQWGjY9nF
3qLk/RY2FiKXnEkFvJcI9+BhtW7Rdz+5kLoSgr7saSJAVtJQQqHObt7EdHsZdEI8Nupj69NYDCct
OHtCnMwUOPVuJduizIE5y+SOGFCqgKAjsjbjdY2qqxjPB8BSQBhQqDp1n38E7kN2Ax1P/B7IFu3G
D8750sgFxMN4cxJsqv7qIq5KetOmhvt9niK3JmB/lZpRZduhb6AWHl3Iyuy1BzF1OYFsx7NnaQaC
V9QEy9xVc6KwdO5A5qMQhSB30d1BYMFZtd/irtDDYDcC8+DZYpb69h9bcdewkwR8fVWhtkenMJ93
8Y4uwl1jHOnK3U43fEW2S4BGiIggccD/MyFnTi5AxdvOXDObFnnsuw76Dwr6FZxNg3VWIIbUBwXj
Myz8FjDjfJBIb/JACppgHBIV5U6UA1BHNiryE4t0YzJytAFiHVC8SopiPBCsYhZ+UfPGCRfKQh+I
NgConPvizo918HiwuI7vMQIqI9uDtinhcaUiEVXUhFPZmUBhmam6NrT+MZdNu7XE9tY/PfK+kdk1
p7gpxrQON/mxxjR4x18KvOb6h1NvWxKyN4BX5xjbNMgMgYH8MC+Zn0v9AFfSY1xgDc3a/DahUPww
5Dktxgt13O8FvL1oqQKmzxJeuHEJpBfKIpdIiU2/UEuqgVE+obDhcQgf6KtDnUrFv9/qrIAOcT85
nwZugk3iB/Hm6YGY6ukkRJwzZg5Pm8a6hrxY/63nvgXJ3eyxl5fZ+CyhGzusF7jgSsQA/KkDuXD2
4l+xA+yOewa75H5Bv8PqTFrwHF58ZFE5frc4tTQ9RBxzskVQgzD77Vq2itx9H7qSVOk2jtlvS+2v
dQ64oPJMmYYgWIIp9aoi5TX1NYH8Jhg3UMpkxGz9tt9Zqni9v1FcbJqjD4jtzk97rQ8N0iSJ2XbY
0mWgb2DtMpqvWgHlSEkxQrPn32EBa9K/FXsn8Qk9jLnLNmONdFcDOldYmbFi127IHw/DvlJNtwM9
fG2Tybym9g6e8d80il4JNqyXrZUJQIhQ7REGRR7Vrcrq99Pd67psVVWBsrwH5CdXRpvt++l9YaXB
Dl8fuwzv2gGJsDxXp4ren4SDBCdnjcujNrj6fF/5tD1BIhUeChylWCnqh0gAPKjsM9lwADJ6di6S
xCLz50Vq/CibbuTGsfdko82T8y/1wzObEyXfBxWeASJ2QfThefEYTHwnbH4wiQlB1sahW3lCRXlz
nUWbCp3RP4vdZkZyAWLs608NhEGQfKrNTxh4MkU2Tf/yomeU2JQ5HPbdh2OIOmWRpjgC2F0MxIe4
4Ub0HRLm9IpUXwrsCIT5mPQn/S8vZs/CgLp1tGuCOEICjAuuAZRNUzidFjEnlbDOPccInRpyxm/p
VXT5X/U6csenpQViNgtmDNRXBDwFPIcqZeULYxBA2WqK9Fg98FPC8VDULvAnYDi1lttwG+sIUv/P
wo3GfJUHYQyIRu4JB2uAAdQ42YP+/97lZNA/OgpzBHy9Mds+ZXrRs4mFqzKPZ8wq5c5hOE4bWxGh
GMXjQpWi8Vsp46QiyHGOjFM76FphALRpaNnARFBhQ2ikhDukgrBMB/VSo4AJzfRBl8FIvkl10qiS
430CRlKOJNeXdgibQH3Eq8ArkYx1PzKffY6gMGu0TwbG3oousNdCIfjtigdfuWKr3EcsVXkIIh9c
K4Rv6hPCw1dCB6DsV+MDt+KpZeZvvu7U5tXslr+ikrDklzm/GzPo53XaDRsn2z4ogMXRJAOYalJU
8Pg0E1+a/2B2PpqrpWLpIReWCWEO97pFA9YBRSd1hqlaA5pM2F38OArQAxdXLrFjWyUAG7+dIA0i
j0RJSyKFmpCWUWm2rCxUs6vnSaxQYor0EapIrM7l/FJCe8HJPENity3YiGTvIVzu2xWuxPu7HRPf
PHtTz5A4ExmkV2pwtNFx+wWD/rp/FyAX2eZKzudWTeWbNtXH/1lcqk2DPoi6fYzquB2mIYpbaKVP
mDpZDSUD1Xkwj6vVob8IidZIS3gjPZ7N8c/FUhG9ijvOOsmVsaDr4XvXsGtTrGPhwpXMrp2GYO6d
l1H8PfzojSeqEUVuk09qf5cOzlbip4Npx520X937fa8PCOwR1Zzq3mBZsnb9LvmGaloL+VOE9nOf
70AeEoo2/vweIgm2m/zL/OYOVQAgzsqpigPbRKZCJTLSK+3boqwiLnJrdufj+5tiSWhQwa34AWDR
BJwOSC+w5B2rabQenN/HLDzLzOAhjOuEkpx0rLNTkIHkT1IJE3LnOTPKfnwfYOab9dym/ILmP6F0
KxCImXnxZVD95yVqAyl2wdZDjxeS483QswqiCzaajqKvH+SdKWTZkEbvElIFuMpb0L4PL53b1pKq
20CduHGCNr/TVA2wWNSxMpicgDqYo9OTPQq/eRksqidsPYr35Op/OrWWZQna7VlNarVlbg5a8qNP
pOcTYlqgTep308iQsyNvv5R2/Jf6/omYtX4w9O9o22sAx91dOVm92ZeAumy2sHJpxC+Q56LtSvlT
1q93wnEQVeEUaEkM0gXL05Z7Q1XLhJkw7qyngzyUHTWIYvSXACCj8o9PlBPyZYpSFuMYIiQdKYvG
I7unm8uyr8ihIUQb1xE5GHyq4pO7VMUdKC/D+dK5Q3Z5j/8GDa40l938eyzRTlcQsFVwOkNUzdLn
kyashHQ73Zt899dkV5XEqjrSwLLeevpL8eZGPO2dJh2HMJvd56oX9dw4uiEXiS6AbxGrV3boxq2f
QFOGbWlZ4jM6aYT9OYBW9u7tsUSH3jl66GPdWAG9PziLcF5wVM/3RVHIgXGhMSz+hSRxBhlu6OEX
K1p/jlE0aYT57bW5+tekhfPJ1vzHbZQrn0NjL6hYFcpb43ww08T0VnlxNhAtf0LbleNTCGm38JVo
1gvIZZ7SzLccl9kDh61U/s0J2e/aj3zDrf4tS0nLtBanTcbsIHFYq7x8umBZz0dwCNvWVZDPMDbV
oG298Dn4S08IlUslTNu4TveqIMCJ00/SSl4jcnpGpnOU1q23ZydNmM5M8xDK3CsdQOs5GQ68jput
LMvJJ/uVHMTCysJ6yhwzUqBs2C+0JSEeNuEccJ3Mo/mEBlmohxfjJaX1Cyh+e1URMOu5T8bWeDn+
39dC5hrbcXf5lKcN5jkS2wiQ4uZXQP6pE6GONu9hw2zNjDt2qUYZcZ6Y4tC0pqKE7qJFP5DALucT
1j8jdNtqM2tU1Z3oiyOIvGapAGsxK+dyhcO5BopvLiZtU5cjsLz/aikvXTWVlc45IrhDTD3A/lZy
Aie4p74BEFO/rNaOeKJRM7VvgKToFIonmEvb7q0lrInnL1bUq0pO2DSbdRApRokdnrS3QlqFLCWa
3yqo4Chtlak8wZHSufthZU/MPkTAfSDCwfmIkLTG3y0XrgZTON9WhHinw2KP3nsBQGkDCNFuT/UM
kQd+NmCPzU/iAD8OijhtmAE/gUiCF9czbLRpSeBZdS2IQ0nfoGTsrFuSRdMV86a2SasKTsWmEiXf
bFFbcYqsA0T8Y4iUagAY0jZwF6QhMAFYjNU7PwQDF0Oq44sENdwfjv11kqj+GEUb1GRLnUwo2dE7
Umxsbb2PBxmm1aVDDi7jZ+mMVgJNxbxFMs3JYv7Bx8uiQU0gQ4pV1cdlxkhZ/Vo6zcZoQlzwXrDh
4Cw4j2g55X4Lwp/OY9nwJ8cJx0yEmSdqBGRe3mmUinGBQJNjBGMQY/gaCvHT270q+qnASeoVsYy0
jC3yihXsL0OK+zJ/xbuEYU8XjqoeBA3L846zyvXeldRljO9Uw08SPKi7lX+uJYUngTNfiIjgdud9
uLneuzL0p55HL9xCxe/ZdiNl2e9T7tdPBi8De2L359vPtlyBVch56eaTk3BoMWugr8V0Q+A4dB2T
e5r0FYZL52kvTS/HWFP31rW2OOVt8UdZqElSyEUiw8cjkFnDTF/mRY5nKlU4+XjyxZA3+8gUnKVF
nmNGkDxVJlF14/NirEVgr3PnQVTQdqUQw/At9IJouWl3OWVlXjKxaPh8EbtcX75LnptLQA5TMbjI
bT5TiQpvnO/OHi2gvgxg7VVxXjQ1FXDfiIPnQHZhqpaFesCFYdYvUScGDHhmsUOoyCG7EsdpG5QC
CsyQqtZYogdEK1tP652IeETusJLwfIiTYDSXWI1vKSvvARDDFtdAbQoS+ud7nvZPhdYuHudYibeB
kcONfZPa5T0PVRTO0EHGC+rN8+2Sd+Ssp0IY3TZTelU6QsQwtnRVIIrYKMqQdvgWrIl9VQjklA/k
M6nEpV2DA1fUznakEUzPrpdbKoQfTwDuerCadswafR6qGLWUUV0e5cmjivQQtBOXUfd/1bzWiTYJ
Cn6hpqVv+O19RBTufw/vO/9FGwSvyMp5m1FdVbkunEamb+lCJIshtf1jv841IzKR5g1dcXNPGWbw
MmopN6wT2UmmfRhJxKd48dJF0NaPZ91dFTGqlku7AuEleXtjLKTEvvnXOEgpYOn1sJVyDMUSsWB0
G8ieT7gIUtrMCOA0OSMd+WM8rzWyzaa2XCuGEkPzwcBkfn9CMSzxU/G6uivqfGIXgBSFJvOvUBrH
svhZ7RtCQRMQ/mLlidXwuIEyUegu6PSZIoVCJLvxhNFDfPZm5oN8YQv7a+eyFHB7vxLXb78owv0E
4iByKi19HljxCNkd4kGvGKbDZJJ607FOtDuJX+TkFfEWkyo/VPCiZ83k+EV8wK0xTuKld3UQ4xsx
5ruqbJyhXKhfD+H4bvO0XAnD7hcnb95FwHVK3eqyxQe/420H6RcoQvrpZF4jgLWgmhuzfrtbWaK5
R1fK07iWB8sOxvCnOzxJyjv44p41wfZTm5GteDUlfjSGAwBDOUEoqYT1ch/Ny+UBWnrVKH+HZtXM
XDdPZs2swoURvPCehUDGp6cqpHM/WPvDxvXtAhH6ZsSgmAVBv0/I5DqYg3LOau55nUtYDhrVp04g
NqCmbk9B8fQnRIBcbWfdGoHNF8jcugVoAwW5yMRBOxrJMxGaTaxRW29RCBIGHoTeQ7V6ZmMHh3Ba
M2no/5izw1ll7gJMCD/IK5mwOPCsoD6Jz1/Ze2WdSGsELDlBfkyDEFOmDOul8wlJSrWAxz2So5II
x6AsSEBNdf86IkoxJ6swtDs3BE5htdbBx2j/cfrYFRhN2wt1iy2CPtxbGelCIwOzobVbGYwaxvpk
p9MqytNiSXFazpVczjVC+guSkXmcRhS9sBmbYVk9mlp0mHMmjDN1u5p0HXB8PR24zR6MWDRmApXq
csp1P480hf58UkaT53sAavL/r4+0++wbbRVWEWnUG27+L9Ss5mQWows9ozOWf0hwdoDjW1/zIs0A
J0ISl33VNBSicwftGt6rwDV6tg2muIi2la+bKPl2w4w1e5/mmSrSsMkx4yJlYI0TfsCitIbUwHhR
z275/3E/CIOfQTA6twHrbGTgYuT6A8hiTB93ESdRqAX4Ijlk/neWdO/b1H+1Co9wrL0nlaTAGhVz
nbm0Z87KNlKNNosU2uI6OKbvxuf0KyhRTImE9cSIzNWA78P/mb46o3/ApUjKn2+6M2Wszmr0Mf5N
yqlMgf7owsMCv6zAlm+IJmUpVi05gJKXVh1oFXjd23ab3laaV07BFv3i5zRSbtVX2qDxZ2EW8Vyx
/8loFQSn5lQykloxCsI/OdF31XK1qR4VPgd235L7xdLg9sII9YTl+3Qmbv32n8WvbUQyzIvALh1V
f6xUCTSIwU6kF7cXS0CBqc3NPf4o9SnTJ/JL2pJr0ufqrQNGRXwZy+nlNRe9q2IeYpIQOVtPiAiS
I270Utov0nMaH/cyV2I95rW7jfStvN8ts+cMJay8uOdLajYivOtmmkUHN11ZSZXs1m1LtNdoFTHg
y0tw67mwwYNR2RdxOcNFatwvhxsJf5hABtVtGD/6OCHpJLNIe8sPe5oUaagIYOvrOG1OKCgRQzBe
8CsTLzqlu21xkwRSjP+Gh1t7D2lwsIVy+pvUMu5TzwGI8qqo+m1y5riS5kEtO9YxV3+510Ri761p
nPNwlMTWZ0WANRtUIBozmh7OXNGc/vTPzsskC+gNDRlNuRH9gKK417wcw6g7OmfUnm3Mp5OKJNY5
68KLWi75NCalHrqjVbZRU+UKjx4S9pxE39Mc8wbPZZii0xF8ibJMyIgGCDlWLT8wbewdnEYg09i1
b/Jhyr4RfpBFFfmoGN8h2NP+xOXRzwdGYUzBMNnrTsXEPfWwM73evHzyJ9Hl/LqkkrQlHukD0tfv
Q/FAOyY4y20VUV9IlKcgObxJPw7OsyrzJPIPkaM9pHKcx81RSC6yKej0kkPxZpCUk+KO59yHWMEM
uLLXKladcb5tHTyGWrULaxduS7f/3HZho0Ceq1nTzw4BC3YlMyVXNu49x+nHkjsZTCCj47oChEcI
snOX66x613KOaotkhyyGNlJ4f1TrGkbZxds14fOmMHFtscQVBT0PWIW+WYRY2SnaqqrlIKj/ZDMf
LA5+f7oMDcVAEdTWiPNWN/ystycUaDcBZ0KbZHFUkW7MGFCkHBY1AYRt/AM3+cPgXPHaqiX0zeEE
wWdNcCQkb4QswqGpGoEj5IYISYAUERwZ8HKUOjQ/zBF69rwgHtd25hWx1bw0KCbMh74BOnFXJTmj
4MwMgZuJu9xsn24pRsSV9KIWCUrWiPVtJl60/NNmE0oX350UMCq8j4AOlW4aBPm8faIimhFgIBKU
EYyB+OpPGaytbitcH1CQ4aLji061UJbM/N0O/tK0RT0n8icZ1r+T1sw1pdER8Y1wfVUVQKxzUDip
Y2ZGGTkMZUDnf1d8dKKEjmpxgPJxiahoPy0KKvn3XpTYX8L9kTYT2M1ZHePGwfHIFpg3YnABqLwK
V+T+O5vrnSgwW2wOx3/N/QPMDQgoJ7C8BjrQ4g+o8YvqeRnSCBZdW2CqkI8zrD2g4+r/KnLpx9BV
qmKXt2aROUxwBPg5fDo/4MfZxiVsXLzySLP6gTLlA0+yk5QFBvPpDdnRJGBOoggLFGjocqCXEpfm
Xko1rZxYtD9z8SA1xnuWGsYV3rEsUTVWPYIVwJMxNi4rWb1m0LMcWmwMdCPjQ45Eipr7yf6vKyDR
Veu5KgN3Krve+WVc3FGK9LHMh9C5WAlevSqDDWRAej0N48ywWTkyf/8MzTTevmwbzqDMOI4420O+
02coOYsBQYN1b0aVqYHihqiYKC7nN4pJRm7OWirYA2YbBu7FWu6sW6drMCo7Y3hUXjIohugrvwp4
bxuNDKEdVZtAdbiM95SPaDl4InCKdl1uW591DCVjSSyAPeC+SzhXDBxpTuIeyB2kdhgBTVHGwssk
ZlSgwOP8PJ6gQY3H/wa3a6KX++c7B/J1PEAQ/Jl0/wmh9A6atbgcaiPhpjqAo7Jm9uWPgS+UVJ0W
botraNNIi2WQnx7Xey9GT4QcP9oPlXIRKvYHHtBnrxG3404htNZCENEOSYxvXJM8W5r9MCi+wD+0
EA5qVZgaimN6HkmFBZvH3YMJnH8EHDkrc2lPAKVcfuRTQQ2GLC1/YEDAHSpbQbguGzbw8AqD8luO
bLW+QaUHecqUNt2m3J4yyUa6Z42G2aSgiytV6h6Aois2yPGhjFK8hrVD7ovbcDBCWIqUC+Hj5K8u
FyxNJH4prfoiXLpd9SQH870Bk3bm/0m0QNLQUtWl9CEzbYNjtxMIMhN1x1Qy9ncOUs9N7d7xARCa
EzJSoghe3/EgFiV9xq3JHDwzsck6vATvQFG8MDuhx6ZhL4zvPQEVK89yKy4yDIe+NvHEKQU5TOXZ
fLZcynRk6RsS19Fdb0YaHGXGz8c8gy8gaLOSp4SE2nHHEITWGISKilPN2lhMcdEdoTn7YMPS7vTX
qqhDlGTsDGlygxgpOA9FSC9zDRLChFzci31VAL6mbjF1MJyJ244lUW4G4i4ajwV++QmPBPlZGqlS
W3E96zXeBD96IGx6FCdAGmwIpOIrMKA08LEXMj/bFKtju7WiK/MPZrIzqxg46bXiWQKycNbhzwfG
PV0tCdDc4I3bXDNUjmTelX2q6f29du9fengFDBOuAw/FehThjMIlF0GuGylghAtBNuzzqCJluaXk
8W164f+FdElWjhswlhSC/5GEh38hD0heKXA4GKky6y3J6WtGUI0qtaeIqt55LhL0rczXkhYF/qYo
g912wbl9RZSdNGnfCBCJNsXYvo7wLjpNgIqJmq/BxahRejoAovBcaDgvkE0TZtvgnQee4SAe36Il
HmCkWb0YSIkd7lUnqT4ZvNXdoqWmq3Y8cHbBhZtOATbELAzx8/1HzKl38bUIaIqh8DRuh1Edzz9a
ojnYPiDwvoXHslUn3qj5CnuYux1sb/Tyjuvde859rG0bxnDEvYT63miaT03utKsg5JRBXQPWcyy2
IDEeElWoi+kqSis1vTwuxO6Y1FaxcIkOHmYoBAJ15vDPqK9nnfxVnrl8aModO+e9ahfuf5JwBWM/
y2Y0CM1Lh+1eHd8alpPBCMygYyt/+jQ9jf/GwqYheQmn0CFWGsxQwao7PBev/tcF4caBpwJRwfJk
i0EB5qazeLYJvpAIKqpusaUNMwP9WcOsCOKWJX4gVQpZA0TyEUjXRKdUvn/9YwnRXTDJYmB38lSd
6qkMaLuKa1bNazqV/Gxy74UQKK8k5+ij8I7UQs2MT+bFriRwGjs4oEZ41mUpk6HnT8fItXAGfwJ+
C4KAoz9+E14t0CBAVeH4j8eJhyAlUkuttfx7Lr2UNpuL0uG2H0L1J/05p5WviONfO42gYHGAK2yj
C25U2C/9zISvPoWcRNrmyQvfSUuTu7lOAkv/2oXTj4kOo7JV5p3+rIktCrW5VGGVXGoXp+uQUrS4
+6Q8BGJQhgq4xtCcwB93SZuwEcR4kjjCYZ/FuE6xltntlNIlmrUAvyeiEcp6YHyda9xfqusyszH0
0n2NkN2Y09wa0EOBf3G7LkXmQ9SpOtRi1YhzD05cpq1tVNQEhfU2J6Gs0q4wDpBVWN5O15jYNakT
YpiR075b/U6omVAZmGgf/lqNMyNRN222EpsemAr8YRvUkzpGiuPTV97YRE5iPK2lATaxg3LAm7lK
rUW0qqqnW0r4EKwCJYruwRG1iqqwX9kryVV+BHBaT7M30lrJHkpj8BHpp8O2wvqtMeJ2/8Dw8Z9i
n0pK79bBscPQrANzYBATeHcsc1w2blB8TZHn9jFv+qhVp/xmj/MMZbsp8JFzG/CKVHu9q6fSAbD4
Y9WCqaw42OCpFk2/3G7bwCl9xT10l4rzui09zkboQ5WZSD1SPiFu0GcSR/9wASL9gttIAxc5awtw
gxvn1S/I8h7uqM5C8rEobXqOGxKc7r4MmaS2LGaGfj1nT+WHp2Kpoh55Thy5gkyP2lf4c/A8uv32
Vbb7cN8WwMKZWJDs4iuC2DX5UtKxGVxDRLGg9DlMNCOmYxzjM+D00TIwAjSNtGQ+tZi2Pja/15cK
+9XagFsB5zQmFhjAEaULNECyf994XX+7CjwdVw4yFKACYnlt8s12qHhrC9376X0Vs1cjd9lOvcEh
/PogSgHM/F7lNbbhKyvuOOzJw+NFa7zLVqwM9Fg6XFYTiTQ78EsoGZlph3k2KlqmBOHhNLgX8QGV
NXMrCSo3eZEO2H1NtBuRSnDQEdbSfcoxZiLxY0yUsys5XrOyA9tPM/L6uoyNk1T1w1OAiSo2vims
LNbabLrsv4d2tppJOI7v98/HrDnJiXkfb+3nqXC9CelLbqunvmJUej17OgfjR9yTHp0T9vK4aKHm
VPDdrTfY7lfFmnjqQfzyvF1CjYtw8kTLnHjw5Vx8A6yU1uW1f3iwUB2Q3y8gptRUry8eMtE/3fqx
7Uj7Wo1S+Gs69ZDWT9Yqb/T0Kdsktw4ZAd60jVVeZuw3stPO7sl4SaQagUWLDV3kS6Zh5QFEv8o4
nMf0ijBV6PRebzq9v6yenNp6zt2PwQYDuAq2cDiQ60QMZvI/XZHv8snh8rvqiYi/BYTPOcgN/wz0
8BgpGANiF71K7k9qgMz8T6duUee2BPSQBDOyE9gK1xHH0xIKsIkH8of1PS9RszHOOY4oikJJiA8h
Q4adBe2tttZ3qI4QDRC4CPMAu+p3FkmMeaYQ+nFd1LQfkj8MzLNWN4GMmQcnf/ka7tNa+aWe3YI8
DFtVKKoHXjHjFB3J5eAs7wqVHq4J4CHB+U2H7rEiq6VSTHL3b5xbvkkX6DsS1liieFO6YOqKRsjD
YGovhhndX7jBwaB+NkI1Z473RPS076eV2xgrWFZjUGx5kgq8Ct6lGEZVmiwYUmWHFXH7YdJ8pJf7
/ImRdyyMCqNLibUNCiZdEtBKa+PFLpHDla5YpkCVgEjhtvvy0yL/9DxlLSoDmFQWa6hWP6vfhZ6O
NeUA70TVe+g8jO1jJsbjqd4HggjOKcu3NvNGR8SZPNtipWhdXSqPyDhmT2Z70YqQPuLcBaNqQYpc
BCDAbrnDst1RCKdOeNVme2jLVuOFmUL9p0BvbSVwTJMkSfPvW7iy9v+nCduNGCMl85frDhzKN5Qq
cVPKbqhHw/qnEdAPCyKoQOF1ASyiUEEcFxDT8CdRu3pD9s1eEy1QyNyKcRjbZ5iUPnFswK/lw6FZ
2/1fI+GVyBd5bvbqQTLAiWCe4lLN6kcyfRAjcPavj+B0tO7gQN8iotHTJWnh7GF6Ns/x+O13VXux
QsGNZJ6d+DjTv1XIjl5ALpfrnVKSiLRqqC7qOxU7wSHqfAVjkpFH2bIiJWFHJCb92fM6FitrfiaZ
A5bk9lOOFc6qc6rYuQW5LYWk1gdyTLYoUd11yilsuPu55MbMjA7fh3vaDQfqPZB3N3vr5+mS9vQA
3V8li5zUYFKV+MtzwPM/rCtgJh4uin2OBc3R4CeH7iDEz9nYLRzccNHUUl/vDgYPb5+CQUF00Tm5
RIJtj0h0Rtdv71tICQFnuNnNuffCY+oMr+SzQJMi7rul1hwpoPVdQxl9I1bo1JOO4EC+CKchnGvs
uIkMync5W/SsFkojuOVel0bin8Z1E0y/uyDW0rAa1AiGfYdfUwRxutzwxDi0o4rK0B+YWTuZRfGz
wrJX9vBOW0hOD3q2O4a0xDJvz+oZga10A7BM3qospQfvKSz+IqlBZ4Klb8Vd0PpVUEIm1APVan7H
hYnBjlCEVYx/wNfyp4TIkYfCQ79TNy6xyNL7h5030RRy/C/Nn3CSqiZSj6/cCRvLfmuEUUNtmFn2
fUSo+N5zPls3GVScpj5GH915EMkr2Y63x/TABknyHsox2oqmKJXtiy7V1BHAzBc8W5HlsCQ4XrOP
raKWJaLEaKmY2DA+KL90wKzNQ+q075wUmMW5Vgjh2gMQMWqKKMlo7EOKf5uNbaZe0qnqc3HIRaJj
2VT8qcZabLHtCgy7V/cWS4WiR68nKOMtwQvJ9loC7j8FOk9zQpbZrxM+qKuTmbDrdkmlaoYdgQXL
A4z96TcLnpmlrPpXh0fs2R34+XhtrO6IJ+znqORn1QQHlcqs1BeUTIeU+lppzs5TmnicnAt98vfF
U3N+9tUmwmmcp1pqV8aQTo7mkF5EU6g6J5I0ZSxqvdN6XQ1+puVnSiDH862G+HTeO01fkSjY0bY1
jV/jrXHCwyo994hX38yIv3gtHOI6CqDINW24cuq86QkwNYQ9mjzMrJlsiRpMbWGJ+NsDQvs06x5Q
VDY0+8KNBfMMORSvCGKLCWQkBLHa76OXvCt008A6YuJxBX652zHRuVaVIuN8i5csw7iwXfW/bLXP
nb5YFDJvK+UNISos7inlNoLV5I0m/F6B3sLrnAUkVadTINWwGMBN2zzX2aCvxmklgllmY5BicWog
DEg+QafY3dlAgA7cfmCdLNmRDmnq1RGUf2Ag5Fn9hofaIt7OJGtRoYcVXnF0pM4bIJkF3mJKXvV7
aDjWs68xSVicSSSiXSR1fBTGXLwa/tmgPrVvZQF4ZBxD2YmH8c6RDau8sWsJev5D674ke4xpMh6r
oCAN0m4KmHIHfCxvWDgC/tWR4IgfW4o7RG2DNvam15b5CkRi9aFD5VEHrBxajcY0WjhDCUD0Cjyy
3sTZMde4wS4D+4NovSWuCe/j6latbjLGX5ZTkENPYSaL5Pn1uFbDJ9ze7qCSXSFVTUe4tvveCes8
0wfDiUnF/fRYboJ+Gi0r/s9V3VPWQZzd9PKZvz7VduYe/jaK3jHhDDI11IF8sZNgUc+1T8nxgIKX
iRpVbC8q7auY326FEuTd2tS3/I37bOwc1WK6PbPIcyGyXZTX8pBXvxbqEqgEzAky1opvjrFK9wik
k/PoI0UhJiMpuxuvcd/UJgII3DaBbXQ2/modXVdbO9yf/IjxlVGApAzqzPT5luQ+fNziNzBZOUlS
hE5ilRFTsLPrS8tps6+H/1x5PfILVJHphPefyj1UQc5eUBHJcKDLR7icv1XfEW4IhmBlXCTUrX7j
Ctvzri8nyXhP/R24j6VTd/qcYAKfUVw1PdB11CltsCupKzZwCMnPDd0eVfjmDLmcDZEdJITlYvnh
scOH1yeUwTYM5+INLUaDVur4r/a9vFeHFPms1550SHgkzZjI7LNbXFOVOsRatD7YGeTGLMc28rc3
hV4TUKkrWZuKZSsYNg9BNINh/VcrHDOPIT6AlVESZqaXM0cM8cM5QUqoElaYKZ7jWpNANHwL/hS/
xUegc7npEjuoSadG90M2qnLR1R0G+d25d3pMKxSQVMoMlyQr7G7ZQgtf9zb40xHeI4VcF/Rb/TyU
hJpkL8bz5IMkw9aqrduqB+flL6P+ux8KY26y6+Nk+nyOnxKt0g1T+Gnz1koSCF4zedTafyr5nSUF
5qF8sFXKWe6vRU1Lwqn6TuZ1PioH/stY1XTac9fnPOfgXtk2DpETwKwPvLYcg9lSzjty8qMTZxt4
azGptpe8eOMTjqlrze5p0j9jFORgRP7QNUUvCwP0Pe0vuGRp6P4KD9OOvb/Z8TLBumtAHM3Ed/UC
LXuqn59zCtaNCFt0AMJsMjrEszlvGFK6eKiw3HQb7LZ/k4f7u7d1/J0CnLt0xULduwxwBDH5+eM6
O/RGojjWV9nkHU8cZu00IQbxxaKIKO1gO+cCS5Av7qrX5UJwx3fY4k6rGra4m2Yrmj6jnwNjncAf
ugbubbicGmmO6KR4ywEH3GXDUxQVluUmMYukY3S9nhOBXg62MdUoXFKPVYbLby1S+P9c9yzGs9M4
qI+xfAmJ8WMB0hrBA2SOy1XTD4ESWk32b9+RaWk8jtNKB80WhMZOjzXw0M5F/8yK2tMJH12GLhLb
fNTRCsQjtjTe2wlFuj059Cn6S7RHtFZ7a1JRW7IXBKiAV74lnA09/isW2SOfx5keAb9gvLsjVvy+
CSFThS5uImyGxcHdrfG28y1ZwxDEWrL8wyfJaPu0AWq/4UXdqwIohQP+uKJi7IYiHAGjN8OiIf0W
duOuH5fXXEo7cF0hbGQb0IGmAY1xa7gtnA4D6CIpilU2XHojNxlCC229TdrQUY+a/guSxU9sBORF
IFKvoeFCQAaioiURBvpiBdrihT2doUvt3h67/yWXFu5o1qlkKCBcs9p5DokbJqQEbyBF213soWPu
xV1CUBpJ0jjtgWZBH2yzJWOBFhe8K4pFiQbIFlFSIbdWMLEGwEJwNBwfYcmM84MN4yAYWFkv2hAH
QZ/hFEPFstz6D3S7hVRA1xgJNHqooDuthI4VvdCROH1HDDXBUaRb1w0V5zMPn79dgKwIRxOC0jGU
8W0fWBdReweKzouaBpvwTf5ZATE/o38vPqctJ5ExNkpmKwJrodvEHszyyukDCFhxDB97R2m3ekq2
GRM/A39diGDy2Q8kQUTNMiYdXh8Lmy0K7x9Wrf0jZVIGWbRQIqmM3VK/tX8tvU/OmyHXGzp9UmPo
vECIM9mBSE8Ni4NtyGtVIyV4St+7ToTY61ITx2EYPDSlThpsM1mQNiAdWSMEhl7jdWCPmT3YQO4h
6Sdfdjl5Uey6632TqaIhQ0NpWnoq/FaqkcpgasWJNzLSjeVckqq0Aqugq1v++1SODE3reXRF1K+5
PvKVA1GHUaT5DJCWfJc8Sc0t/ksbbzSxMj/+sKFp6c5vqXEb4kiU41qJmOa2Ku6nqweD+WjuLqO9
aDNiGiKb29sasILzohMIMnHNgEBWEuesBOLnH7DKxQPGdA9AWauFN/rH2+KrN/aTzjCyKAEZO+uf
EAoZMzX9Fgxb6sHcY3LcwsfIdp2WRZtTTVCMEbLw8hoxABXqLhkHzpVuRnPua8lkuOPhQoAGz+Qf
yinlCIPGr7VaSSO8DxXVppkSt8uBrhQ2I/xlSn2YsrcBfeuYVJqKcz5LzjOFxv0I0g0vkcwQTGD+
UB5z8FN0gJg5qm5Xz6fD6NPiei+J1zOyTtLHB0cVmWmyZK5t0vDGWeFy8YwRXwE+2JD5pa6zsI7z
4xfWkjifNXGOiAoAIuq9OyJ9DbPK74nwC9F19hG9V9qmk3aMyXEgKiTiXlI+hdZEl4it5EsoRVW1
d5j33BoH1k8KwRuLtK1f/aYSNQ7PhzBRIMZBXqbpCbZkCCcK7F/xHSCtAbMNO3h68iy+34iHsRd7
RzY/x5tfnrU04GNuxBrM93ew8OvA332VJE+Y0YlE9DR6cOeS+Y67FDpS3tkUkXj0boq+OfcQV70g
ydec92zC6slcHVdMKdLiM2K0h1YdpQtGRgszupL15gcLJIYkpwAo5gBU3/POwXzuO8sU2QUw+sBL
yMDaRr5ALgiEmUTIiCd/WkrqgqWao65cNJLJhp6SIfFjSxSLpvfhzSCKj3ejOBALDHz08auHUWgS
6PFDXflHJDipf7be9km8Qns43gGh7HnAdT5up9peFkbgmm4MDzpNVj93al1MLDY6vLy6APrUKzxV
tT3inkqN5gMGVGxAjV9qQ+cW3fZ9dPFwYyb/0y6Sp646jfrhwFBzV0oChCsC/cQdCmHjtqqrvA7+
ukPtbaeEjPyIoXnuKsox5o89hE50ShjcvAgAxPlc+RG5UZPm1yTBCXAodFIYPqr17hfOm/ajQlhQ
ojB9IqhpUm7q7iA9EY1uJiKH9Xnkt0o8tx3amR7aUQvzOutLr74G8FMvIE5/Nohgtjt4FGcWID2G
iVSDofkK9n+qWLe0z/O36z5m1eCwWyCJyPI2ZAAGqm9b9MYtoR+YqfBdOOC47iHMGD9CYUp2SuYP
MbNZI4Jz4VYTH6p2AGPMx/Q6/bU15Zcz/ID3iu++jE4C4a4vqRijeBryvR8uxBv17sfdz+Rw+67u
LjbojJDoCVjqYVqjcY2IoIM5UcXK3ezbje6hARusaxNva0F3eLAG4o5DbxcYnGO4d/tc7JgtXvqe
j0CcmUsBBF8w4I/e/PB7m2P956aHVRr0/CWX7gPqiytHNEUYJ8HD4rzABE1m8a3yGu4XkM0MUaVm
AsvPCy5LhExzkuES6L0FNjJKGQQpvkk0JG9LpD1pTVeXFzPCpx1yinP5cMwlqm3w61tfIyqNicBO
BEJRdo6o88q6XVzhUrWfpytl2E9Zo5S2MCywAr/aI63DCUIaGe8raswikX5VL1tcMJISPsW9kgx+
rr/QBgICENWFZM/7Zyl05Vi1BfsHVROX7LT9olnnl7ecXsu9MDAiSnxHNF6ALCNjDo2ez3YUfsFy
ad0sT4wia3GpZyQQTQnycw5WaTd7Nhc3dndSMgYfJw7QaNM09DWMuHZd2XUewJJK9IMtlAKRwW4E
1x6uJ+Fc9k8zFLGDKK06niybkWKlUNFCPnJtY6P9HapjLPz7GWdjrqptb0c4H2HfwIpKChLSaGDE
1Bp9pgqkyq5cXonY6YMBwAmqnruRH+8CWGhrZ1nWkL0NldaxaStcL2meoWz5DqI4NHmG8pmTEQOA
3Eb1Yvuhb/Z/GmR8J+bxgy/bto4W0lyiAmIhNo/PJPmgpevvGhDRxSrVTqfPrWjvlWGByEFbNnC7
RS5kKUslzCNk/973ULu3qYScdjFAEB8nN7aZGeSbYuac3+rJQziLpEk3bVhOfs8sJBuBxdgx8/jJ
AuOhTvK1A7Fx67u59xU5nkilakgHKU8f8DdqIf/bYgqo8Ojgv58qnvhGcMDhnnu6Wxstq4T50sVo
kEPIFmZSJzMzgAOYWn9COwt6Gj3gF4PZOfq6ZJOkBr4GZwVOug+Halt370EL3SN5VRWxnla0Ens1
KgBr6/Y+zHcof7+SUAKOP63Qo3ZoJApAaLQ1mh8AUyEwz4uRLitsgWVMyEnFEW/TeH1S0qMuE6iS
LthLaTqOPxpDxAcAjjFi/u83LOYltccLj2RUEp6S9bWY7RxEPrUXsNRXC+XyCviJqg9U0gUEdxBt
LQ4ie/K76hLAV6blZIREDUJ2sINev6wXZr+KsnUp+ApSNPA8llDb9CZAjRokwe8F+KrQaxtN+5vS
JEW5XGAcVlKBAjsDlYcAoTy9pVKdVsQHRkZhZLYyPhZJDZ1TU5k72ksPfsBk0bME2MPc4Le9RJcU
jUaJDNL3qBnXHOvBzrHnxE3uMRTXkLQ/EqWxjrMmuoYYKx6mvXb6PUAL8YqMUGf9k6Dov3g1eWnw
jFlrDn9J0ApKaDdKvMmeWMRm6GEKTQk6jPmsl9pWmAidgW3aab+SY1eYaqtMLCwr8KXb+3iKEjJh
NHW6eo8w8ZhOvRvUGV25kmEE1pr8+FA9Rks5AfGI4guwLTKWIbhEstgvAe4IjkZlSy/uy5uEu5+4
DAnRIZq0Gae6EfEcesDyU6oivEskh5GPN0+U/AxdBsNTZfBA1GLP/Q0FSDyoyiiTt4mF9gWbFNZ0
NQKIHQxvQsrGIBs6EPOiR3xjt/pDYQnxVz45WS33GgVtCEbkzTg6BCYysMzfo/HlwciGrqzJkGXd
9FD4NhvogrhMuTxd0oV76tJEtleLOpGEEOFzLMvpeE+V7RzZ3/7R1Fh1bY4AqYInfGIXPMSlwvPO
V6F9GcYDZ/q9jYeM69ZdWmQ/VqW3zVkQ6AEYam3GvZ0vqesbG6z6HOE5lsgPZfloNeyDf3y+ttyK
PNlqWPUY9uVYDPqEJ22l+cJtGNKaDeeDwwqK1Tljto7ka4LsacPZOn0qZh3gWqCEvzEWtepwpROf
Dc7ZzPkJkNz1Y2KqlRRxhFCe80IEjqdBuPFg5mGNgddYkfEImaVWWVWzEpAdE6OOJRF/aE9+Nr9t
j2AsXRkqt/t2eyQ3N0ZQq1hMU7wZcOzrXTSA8I5XbyQhUN+k/zVVbSUh2Hj4QboYRGurcSnuumQd
JHf6B+N8sMuQ/csEmvX0MQ3QYQfQVBgyoe/n+w49/EMZ0JF3Tgv8pq10ojxDIeQ3KtPpM40LRdGG
4/plM93JHIwRQ7n0wZs6l681sukBc+StxPIk9E1QK0OPZ8/t5HGRmf/b8EoUV31oTS2ZdEWT7Mzs
h2a9QDoJrdPOIKMKFxb+logDirQrR3PBkbDjW1adsrELREbW3IREYKTM4X23c/8LcxvKRM6qjCbd
9OPbke46v3s2x2QtHrQCE8cDLX1S8ZjSb7jhdurtFjWw3slar22TJxW50z1fzMUx0CdQ7vwppXWc
2ibuuMqCX8vbIYngrwj4W0rE5weR4fkSEoVil3dMFiudxPKfpBfcNxlWIMz/2fx94UAo00KbLzGU
HzTYqXO7NLM9X2HNU4HjvEfYm2SIK38zZdNQnojJe7L7uU09evqtHwu1PQV8dvusKARAoCWVy6fA
AfskeImMxJYCJxc8m69y4MFa0XOn6R6BUfwT5LQN1WqxP0Xltjd8bxK85WGmKERTofh6rJD9he0H
AhLBpp7MjctFhTDWuMXKnuNz+dVFv2W6HjTowgrHQfwPWQqm7U/8IHeYTf96ukQV8UB80b+QBus2
32EfgVV914cxy+7ai/qfAsj3AB+cC6XZqS4DJcniaFMG2AUTxDAwWY5F4ppB7Ko5mRBByk+GIPmU
VOlM2z26wmEJKPZsfeQA6pp1J/X7MklzewdSFH2syFD56FyF5SlGsiaV0n6dFM8PKOObRt8kI8QZ
M+FXoFVMGkA75HhcEVK89uSxoXqfmaaS0X1JkXXFNRzVc//KxRjnj/fybFJFYqhOjKkLU6r87iKi
ueIB+YaEU5kn718zVAmV5OyRkRdSdE3dqho9LhoRsjxarjoYsI4DIIOkLlKCO60/P/ed9hWp0sAe
ja4Nh+lHNQxI9gu+2Oc5pqsSWWVQN/GfrKqX1mgZoUfmJ8R6rRHVCtLKfL9PUIYV+JR4LjhWA7TA
iirYhk9vSVEXraXSxuKWDcd2yt3dg8Mae5ItyJgavG+Um2mLa9r37TG6Yl25unSMnx8rsMjihpdG
T6dWvymF3uju0zmtFL2lDAN7Y8U6BfVBMq6fJjVJSpXbW1NdfMh1ieTvBe8fdfnC7KjkvUrZnaBo
pxi6UZLzLK4eNdRdBwtvPBAA6xTr1deRGBPT4Ts+v/Z2E8Uq+Cz9I8YXbU9CYlziUnqx1cLAn1vx
cc2DtJ2PDrSFABfCicjKR4T0DuNc5SOp/ifB8jvXruLXFGhIlP2AD8cCM9Wtvk3WIGYXbnwSA9j6
5ks9F1GRr21X2yqe/f50TIcivT1ZAopamETK7qPRFbaYaVnDj4E0YyQ30qNklUJUM3RPGXTRmEe5
drSko0M7a8FQuJuUPPU21pWKlT8qJzDBn6Hnic8JtE+y7j747nAKIn8TU1J92et/bsh9oSTo4PhQ
nQpuUCErqC6Mn7tqS7fj64qm6xSDLNunSy9ywCeSxTwaRlnjqIOuMbNCypaDCS85oSQxPQQh6/EA
Tp9kFwWEqirfjdvdVM4N2uoVWLM3Ku5RfDGkigj/1RWR/QRBtYZlYMAcXrtj17bRpsECEMs+wS63
7kbs8m6cDfBCo2HU3xDe/fbqTqEm7o9usX/XjV0mfmFnD5/O7GIlGttm3MbZ4kkQI0WqapsOdABo
Z55JWQMV7Iah/SFEe9Q/Hd9ddyjsLyQUNQggi6/omzEtnUNdlLAvaj06x2CKGjjeyTQV1O9cE92T
xGyYGdDu1TOvMBmHpTYAiaEBdqN0Z85mA4mT5zqJED2tGrw+hYkyF4pRXoJjDe1+PmXpllLBfXYG
mMprvT7gxIdiMT3SWsr779Jk28HKzzznJAUye05gKrEt65Ufa77Uv+AzbKV4niXyRDFp3LE7X+jM
DKAwAvp8aMBxZFFes4WUqmkaVL4/WeGA2tIraQ20hwtiY9Xz7DNt58EqhCTJ9WTBe7WyITNFgQms
4JrNoXcpgQ1T7zzHanNf7sdLv2vXeh31eBt31JGDh43/Qk+2zh0W442jlekVBKMiCFqZSuTXDeQp
h+mkS6CzSJs9evdMhvT53cZ1Uk+pBhgyjfuALCW80ZTemjXNC+/fo+pWBjsfd3/cRnbS8X2bG8no
g51i6qpIycv2xa+pj4G535ojeOSjVE4hufAQSdtmNReQHeE7uxkkC74OMgmfNNrY5lmAiAxSmK+s
0I0/ICo/cDKy3s+bpEbVaip2/i673Hz9F5sqml1m2pYFdmuF63D+CY8/S0X5PAkmz+YlBzwKBw43
RFhtsxGFG4QS3wehe7OTgLFOqXrhc5dsgpbBqz509H4PSSMvJD/hsbqp1nh7Jy98L824BQJnZttu
s49LTgDgTgusNv1aVEaqYH2oXWuL0XwPHIQJ6tV/gPcVZWEWfXWBh4TFH8r+kmVSKY9ZcCbfsUKV
OO+kQuDuLpTfa5tL0uG6F9n+dn50sTy6/6+QtAuTgnG0bs+OOLvgPzIttQbwSGL0Lv+Caz/kIpIf
vmCVOjpZ1kuOOhVrqBdLIlFxVGBxE1k0g0wS1rZf6kXef+FXt6SfD8xD9vNJQmUK8XFLO1cMOB/V
bnIP/OCy3LcBkPmYNxH1UqvDxx7FrfENQYv9BvPxl/EXOd8V5ZAssVMCqZw9HQYI9EC2ilYc7A1c
3Fp3/TtbeoiZ3FT76S186LNi0ifq/P6vvCZkUmFu2zymCFjYcAt7wWnGn51Uf2nQtjs8EAGwBIZd
4iY2tCqPm2hFhE+GD5LDPZJKUb9nL+P0F7oJjcOkna8JhOy0kNQMZCOp2qqHK4Dwwj7IiOvC6U+U
jA9b4FcJyfVjsen9tC4UyZxHnIJGMcc+LSMTEEaX2lzb7i4OQGwwR2F7a5y9FcSuSc5zTGMdoCZp
+w9ENT/hK+MMGFuc/qowDFcso7mnZZjtlTmpwN16di5nCdtrmDsFd/iJUI1fe9W7fztWgXcbU1Vs
Wi2FhNnqgx8KrXrgOHVKdCg9aC4TpYwCe3nFcnCbSKy6MvwenhBbQiHl3iKpuUkS4tywXuzyjH1/
FgpYFFuQWKk8fiqqczLM1mG4dvS+yOwdqcKFlu7BnnY2we3A2Tjl2HgsfNmeCKzSwqqH/8rKEAP0
BEpaNkvGCTjm1wciGin21edAg+HVLwe7YJDI9yxTUIkIekUoqiws9Jro+YHPVKhEtglMSMEyKvvL
cGpRcRdwZSBjuFG7llXkTOS+ZgQ3ALqTJLQL7uzYif0ktK5b0IHmtquFMADXc/uHU1ZCGbWaMC3n
bOEuxUZiufTlq2laQ57Z35fBy/vOA3tdS1pnXKX46uyZPVQ0iearkOSM9zUMAjrnvRl16Ki8ndzd
0W6XxmNA+LiFzGfN7/LHnLGX9bnuUmrKnloMrzgf4+XinS5FRaLmTPsIyAE54vSbX3aSt1dgpTI1
Jz2NHCX1es5tmPlDWQfRkiyIEV/eV/7t9bpFvo2je7k+JNYbCeOCHSyP15B+2i+7kJ70AGXyhvEB
Z8YqUW8IT+UX/lAh0SLBGLWqL/v/nk/2lxDxBgCYBYiYoiFBuc5fmh+zzJPXbuBurCO+iNtTAUXo
ZbOYNN/ywlYLTnmdV6AtFENfmxhacQ8BOnfX1X+UKSyikXyFo0f7CQsBZQFFUcbVPEM08G2XAEJI
Koutw+QbaEcEyB3J3sH4rRtwG6/HYjE2CjmLj62QC27w8ym73cp07KOn3mtGL6NRaZYl8u7jM55h
l97sPnF356mA2ZDNCYIzV2APzI7ukgRyD3bnVVoU1lpS1hJElol14/8CQf9klRZNCOHinkH4A4ir
POLt7QYnd+HolhNzYR7GoioTEcZjEYRgXRVYI114n+xqR5IFPZLrRZqc0d/KqiexhXlgdtvILchy
m9HXZ7DRikNM+b7dhlFLPSQWvMRqJ/c3hYcNuI4aWHOqNNTxAYRwvXdCOz9nrG1bXBrxJSXfkY9l
eSi/9/gCQhIREC6WTWKoex5DxnR3xYPuMzr19elQqNZyEDlhn6wMZ2ibOWrDvOj8lF75uxlnMq6X
kM79MtrYkDm8Dg/RFicLsPW6vY+Z2My4j9x8+OXbhA8EslpgWojZLLDE14N4/yKtZoE6adizRkie
/ppTVJ5/fhBb8fyMIOC7yILZbTrvtImM9Wf/+lq+Xk5q+aYOhxKs+vTbmj5wDlwQv+KFw6otIueX
av+zO++Co5kOlMgiHVl8OVknYesz/lwvnZNtVRtdlFdMmBsUkMRoAl6ng9k2fsIe3NoH4CQ6/plx
hA3FiX6j2EDnrffgyTkXlOz/ZK/NGcVthtaw17d6cAzjzmV+KIElPLR3QMqN/hx3mKuNFyJoIxxY
D2IzNv+6nnqOs2DHj7tNMwrEyvuzqneiGZkVHsQCJAGle+8DYi3eZ24uLecn5o4rIKmcnywfw+es
eCmroCD2jLpFY7aKe4i/9oyV5UZMP3ltM4aiSX43h4okpRmmDcnbfUUHQhb/jgdKaJ8EhZ1FoE10
gfvwwvhPFI2yvP617xo/XQ6NsBxQuesaFtAmqQ1PVAK7neUP2iP07FZa0BYNXhB65f8QynjMxUXQ
FQRNU4wxyAAhJA3fEtPAPVX3AbbO4cLzDYdLrap9rEZoYSreKVLlSlWulfghKqFDzJrN5H+YSAOL
v6DY9Hfht/8rJTOsJCUfFuRP2KpHikcUF1KkiNOjvRF37yvaHmkb9+TLH2xer8rKHX/acnzZeguR
oM0paoNwEnDIm2nx45Z/rM4rUuAmIp0f2sHIaEQ+hb8JTrrsFcus8ttP9kI6j/IGBeEA2PVPDZg3
aJ1rLwLxsxeYNjOZxVAbJxbfRn6SE2rKAGAz5g68N7D0bwob8Vfcn7UiF1MnmfiUKxiC/vmrnBpQ
jUTk8iqzNzSUBoHEv9EFNTuKZQlPM39rJENo6STq1kV7bKkLgjdbpp83q3oza8/rHIerUfE5yt3s
8Rc+056Pz1R2cZYoJ4pFCpRUwBTXLQR0i0qjNq514Zo+D0GI5ohs4pdz9+QqIXJVnEdk59iD9jqY
i3AL1gs8YATgHXLmifFdeqf4+VPa2sxEjhQGlb/YP0U7PkzHvgW/ilLIJCo0zwxi46u76AuQQwHe
72BEJLoqo9eNPQLKnaM/XiuMaCcovuURabB6jq9CiioZquIpNz1jT1W3JUQx1R9LEttXi3mi49Rx
gadfDPjN/hzVwnVPyf51I785Ze8B2xcwz3nWzQ4Nwa8wKiLCWkwChLrZv2DvWPE+o+kanZ7rsFBH
R30yq4H3R9tzLbvtVzP+5nH7ELvH2yQrFVQo3AlNFII2pBGPWkntj+Rfv/9yx3xRM2HPWijnzVt1
gJxu2I7OrNC/cTggz5S6UDnJNVxUkBpY04+wSPJY4kTuvMXlFnLpyDEcjs9khpo9bM7ixd60Lk6Y
kXOwzs7/vG9KB4gXRPajtXKp8DTVhuwcLQ27XL2rvNngWgfvSsMczkBMv3xzbKHuT0wwiqhNFkDq
1TY+N+WT6ifb5xhXu8rcqZJHfQISUZBh2eI9lfIBHdn+yaBN5ZvIXtmB3tABibb2/cYjwMYHLrPt
Tj8XxHubaV5KzrWiU6uIQCie+0rFpJ3GX+x6CNGwlmq/GyDZOQhGsy8vBxZ4vJb7muq1nnJRsrmY
B5CN1KIaSobd3Oox172h0mqZpZ2zJ1kIuU2R1nUWSRNVxeID+YmoF2Uwf2fpEYiHF8PYd0e3ZNOK
EIobyGuaIbs9YDUZoN/nruROrj86oYamN8o78f7rKlhD04IeY3vkLhkvYyCq/E10DPh+Fn1pyxqb
NSnKh+DO0PHS7ReAZL3/wSNpjUqKD2Ioo0FDtv16ZvuX93gJFpKlC/Msf1mUlxh3awywSr2D/v3a
fM3otgDis+LvFl9ddI+aRWwYBvK0QgoYklk4ZBtCrAwMtnuW8C2jaAz17CeIXuMWfdLPVSSUkaJz
b2CXYeT+mopPx/gZBodmS+vwyQImlNYWlrtCBmjTfvl/FqqGgbeSG0hy1N80Dsmf66pttyU19BXY
Tk72oscqxVIESLAh4lunCEKF8vONoTHUcKlMugFeYQdlqyh5fqgyqKa15P4aQxnmKW8aUDz9LT3e
nNLXlH/yx5o63oKKTixAIezB/dwSIMah0GxpqHswVtfZn6AOSnbf57rXjvx/mnIZtie+0c+k289X
l+CXaimehRW/GMYb6ZH4yqEcYRaKdvu/7RRG6d57P4wGqxt4bbDcbn7j429fkTcBHjeHXI1NFg37
XMOUf6iE5m+SYGm8cnuhGDo5AszrImT9wld9axm1lsWZzj6KnepdWD79H9+0FvkDGpwYZCDMz4F4
li81dE9Fr1tE1Y/4RNQIp/2MUh2vazZT7j+1PzBVWJuYwvZjdXfgOtC9aDysuDXsGb4bHceLFvPW
pU7mRjL3uAW8MU5iJn0Z19bqlT78IxZK40kG0Y30Ub8/THJfONhcSM0rSxIJ0kux023cx7uGXlIM
QY9SdzMTvXc4KNKppl4FUl51Lfiw392/NhRBq+15zhumuC9LCealXLahwl6izuUp9sDHeloYhsW3
sdLhQ/K8DRZFBOHQoqcgH162gLLGj0IPtTYOQVrJscmtF4eDJ7VwRyboIArbSCbQ7ZuXzLltN7xs
Gq46hSqsUrCDjDiKEq6ULlKmqj3Ac/ePSak7be4dOho3zMJzIdKLax4MCahj2L3KCBHhrOJwDTZN
vauTVbnqUJNgKOCefErCHCrKMcSuw+m2rUSEYzQZ0t2ohrOrd+01GBa/P9eQgBzHDkZet8fdx95t
oDR2LKZLiAtDTd+IGgx9Cgvai2vszjgeevPtlyHjzO6jpty7UCAmuF65FP0Tt8M1V1vCLPUXho2/
zmQXS7hkizTK2/0Ro9Zl9z7v0+D/W7K9UvLsjmKsqlsiBmy4uOQHoIyxW6GjKXzw1Ja6AIahXs+s
5nOPOodN77VbC2TVqugLqTIFnouoBgonGCWpgpk1Uf1EkiPNFBp6Xmjom015a5QhNczK/W0bFUeR
mTjVbSjG6UlITQqKjfQjN4aGqdBBpQXfTSlwmU54TRaSZn3oYJBnMe9qiox5QNZwOMwCFw52Do7v
Aslwq+EPLPQONCeQunusEMWWNHHgInlR4+FEyQt/sgrh6hYCtyL9Ixf6wEKCMJh0yt7l0vk5Ftwb
U9I2Dv8QtLrNgqHdpTTYolvvzk7/DW2DIHNNVTbDWFoYg3iGUI8S0ah8fp/EkKwQoBFNU5YhwOeW
2iwx14iuIt4qo6+qWe/7XpiyMXJb5prlWQJOLvDE6O+QC4wvPgG3bevGO7+ga7J0uEXd8YHOZ4EN
2bDhaAh53fjyI5Rw+85funRG/bWtH8H6aJtzFUpei1RxdhmBiMGhI102JBq41tBGLRHwPg6Jw8DQ
EdDdPTS6dobIZf5PACJCsj8YbuNezQcGQGR8ko09o+wxb+jpvtQv0OBJ9IwXSoUbzgJZXJ3qjLio
9mE7gYjb3T81cJ18wHr6imuXkQRZk1WeCGGSNv+KHWqtKKxLEM1TgyG2GEneZ4ZbMl7ne0Tk4Tsw
XjQP6cs8wRZnqkhVtzd3/xTZqdsGrPPDkokM/iN3VDzLAaRWsFQ+6Skbbvd3D5gNLDmTvjIIH9ty
M6l4u/532wnhiN1AQlVtBLxZeREVjI50aeFqqewXJh05rDuhiFthTaCHU71VGzPmAsEAAeh9oKV0
7HO1z2lEDumm1mJTQCqP0Bo2ClDcemGHBnAkbqQGkEml2tyyx52t4BBXJW0xh9bpocMpiiemcvkD
5ZaLUScDE/GW1weH+HU5u1ChP5l2Iwrg9yB6okMtRaSMIfLiGcyukak0rl1VQ08R4QX3eKfRNCBy
KP8f43hlSVkAozatBMk0tgfbTcEPDqvn5tMiVoDa90uGgjGUCe7BGxsMaacnG3bDFjjnoqB9RiOV
kgvjzMDwq2KaEj7xgcCYYsituCtXBPByw9/JHw2v6GfuuBtPKuzrckADlgCdhxAjYBl+p6WdJg2o
RyehGvgtIHLhqjZVjrNqs1VE+a+RFgp2logJ5uUYYUrU8I9UdO3vQ/496vDCdnr8/wi7f9ffBwVj
c6oVuJ0F4H51eDmY8/vIMex7379DjyX8f+8SmCAyJNvt+n7y2a55SweykCKt4+3ImaB6VQbVxb5w
if1xNO4ljrC+WxWJZjsHpLpU/GUs24c0mgdigpG+B/paXkZ7UMK2Q86vca93XZBfSLpzFfl7CRrv
S4+sHI/RzUqIE6QWPBY4aoUtjGbN+50lCZ0TEN97btfYdAPisnnyiZT76yRwxPrIWNglQVmhFM0o
jOpopLLy0ye3Fs490Z0gf5CTFr2DGUTtZ0juO2yLI1Azs4EG1nugzL3XVS8dkwuY8tLVxXB9akIQ
zChVeCJXzbhsRXabG+sxCsN/QCBBzh7JhgVL7ds5JMNn1jUOVXp7/uC71ogAsYEtD5TzDVILbu+L
KJvoJYHRkSXDT3DtJv6+vJimG3Zw0kyxP/f3K48MNp5OeTfzY5QJzBUku44YnxQwUCmkFQG+DBEg
l/ek5Jyn0E1rXblV01YJ60ecbs989iw9zq8uNEZxOAq88F7wL+/N4KxRLRekWAzGQWYT+jrYi/ta
QoUjjl3IDXuFcrNBXzJDE4unWR/xRK49yX92/579UU0Ww2scOHAaf/JRJd3CVmytOJru/ft/oLpV
w2Vb9oYbxxYF4xgrh6KBthHkd1rm+Oc3uAldVzGZBWYorXWYN1+AQmu0+GTBTwBsybR45QWEJLRR
BT7S4ZO/ky2ZQgSTcBdKyz3bQitaF5AMbr3dhhnZGNFZe2JzG5PodhCh+OGkRJj01QOxobf7XKbG
0bNCQrUvKOTlyaGwgwtIrdjwgaXkOnFJKAAu7ONDvTlIA694DbytCOVi+EFvjuum8ove8JXL1xY1
0gnhW1rYRdIJRRSMa0g9lkny+jID5POGF7rIHOpdXs7A5XwHEW3rOpxZ2+cX2Eh2k9eiEDIe99qb
CBVNO3g7Ddnt15VYm4KeGaGqgyZxzT55VVHiblcbxs6yxZ99HNBQP9fqpcWr7UmXhnh6gVxEqj5k
XJPDBzAaXF+5u0Ozu6i8fJshS/hMZOMNkyQ0+z555avw8FSs636P6tCNiWRFCQHH5kG+FxIzgWIQ
9fgVxOQo9xJ3L19BX2U3XOSlnhWdpMWcSAchSKIhEIeYbng7FAjBzf0Yub81ByOuYUAl9GHlFjkf
cfdV0OvHleE4meGIewGtF7UWvSd4OC7SKWVZXHZXtNTvwmsj6pcbfA8aY4w+ydEISKjyX/eTev4q
NhvYSddvyrsAS5+aOxZ95DmhmDTpIin1nZcwfjYMx2PaRmK8l3aEX0oaqxPiPu+YOjNHG1MhFCNT
TzQBjz9SlRaMxWb64qO6sQrnANPVCD/DB9ZmKhW/S18L4evLs/T7TtDHCtOxuclDC5ejRY+cMRmn
xdj4gKR2lXQ8vDuPfw+Ep1zJC83y3sP4XydA3W2vr3qvL4kwZuVv7la1wKRLaVmKJQW9bfe/A+++
vMnHIBV0OWwvQYr8k0a6tllmPoMDScPSTw9c0P1kb7raz/1NxQAgQ9l3VdOueFsSstErFoJ19Wn2
3CbFMhrRc8979DUiJaU4BcofgbhdidcUXLDh/9ulhOfzYGUorBlWySYsM0hjkt/N4kSXlASbyXCQ
XTxkXRJp4lhCrBCs3ukrZ/zTPvZjsRm0darrOmRUErGLOAId4RkoedzyJIeMtWtIctHO/LiK60Lt
NpMPEe1fA8mBD0xVSZjDNz/5oQzXJ3gLOEqRWy9/663GtmEF7LCRX3xIGO9hjBqoY8xjFOW2NhSq
YmtK96S2h0USbTkl2Hmkxu8T57CYKHNxJs1TBMUaGwqBJaQyxVlL/d1nfHD4l68Pxq9agABjLbIR
oLRhMoiWt1JXaep2/958FwGgfiQ90AXmB0PMw6rTlXvrT90xuNagxMRwQLKKo2Y111MLipONBDdX
dqu5CiNAxJiAxF2H8oDAETgOIJKqdno0r1RwvnT6cXPliF3FxpGhEPG7h0SWyeyhk3eOuyqY1Vcw
FnYfxxz3NqSLQ84TiopwOet1u1zMNtx6DSqa9kwjPheXVaav/DEKEvzeNU75d7WB9qIabo2MXVje
x3RsFhE3M03HrPx4zGpr0F/1MX6ZTCZ7/AF8Em7ggd3gi7+nQ/B8JvaB2cWXmhORZVtik07zovG4
XCpSbyg8VJeyRH469eNpGg++kMAVIc/ZjWop6o4Xtiu6DGK6eNpprRhs1csf3Xrae6mK+slhP2q8
e9r/q7aB8t1j54p2IcyzCgSkWXoCdyJuuoPggauCnmw4dpgNESgVmw5suqV9T6yO+HOYuOYFmmLJ
bJTJjvAouMwnL4M8/ttt8xXocC+I2Z71cs+ClUE8OteooJU/iNsXuQa+TQcu8dX79T0jkXIAFaW9
5r/oRVCW28dIBO+gclJPTQGX+2RJzHmpE1r7mZRkg5QquK9QSTYPsHVvlXzkZS6dNh1C/nj6qy+f
K1xYLqpKYHArQiS7w6tceQlLN/A26WN5J60WlghXA/+0Pf4j29laFc2/VD/T+dZnjbUf6v2G675u
WdV2Tis/w89sHIW0UIt7V4ngBX9Uhydc4EMY+JfPLrCTzPxx/1wM3aWOk8f7IcW33unKECFU3BQE
iH/C8jkKE1j6kiufDyc+tdB09QKEMY9oXWFg/metDlZZZ2OkZyolIelFtmmq0DNdXpAiGNiAzjVT
nQWjdsOSmvLbqU6Cx+YfOHCxYttxGligOveR8up/p1l57F76Oy0XUWELrkq5x1kq67NOQ0nZ5p7o
yoDMQLXL9glVwa+0UKFL96co7kAZJ5R2VNaxp3fLtn1B883sWmVFEaXZTMiBCdKF/d24sO2GWZ8Q
x7GghoB7ZNfTuoIG+TM3ErrUkvEGUEteNL9cJoxDoVw9qVpDaWndo+9pCqa6G9AJpNI7eB2Tiu8b
znsNbPnYZWgYyNJ3n/ZHRJe3qjZgP59tbJRq09bCCDqK6tfa5SUXgi9+FJj8SGvP7IddDyLlGNxG
V2OHxg2xovAWSmlXg0n1t9JniGDpWwqEyuxVlqr7sk+x05aT6p20n28KIllJAE1itPLPmLwvhJHa
87dqa7gO1oiDjn7jMthABoKwTfe3lPao/ln3yh+Dhk9OFSowg/ZZN0DvHOUuErwUQjwHlDakr0sI
J7vX7MP/2AZczQLa9SN6gqb3FGm4yotOrJbnQLmfASwdbGfQP96TGRV/aFsZ0hECC8y4fAC+hfkl
00MMmPPkpoOGloanyAO6EcWgujTiauqw/NYb7wZzpFKhdrQ/6ASzYALhAxJVVSwWKY8hl5cJ470l
sXucN6Vo8srzyA7konqimoZu0aq2E/8iNLPY/z8SQFzclX/2r0lGgG8qLXOUGaKDKrFur09bWVBw
muAhLCg4XEk/LpGjFb2ocJWd7Y42xqM/2kYnIogG0UblXmQpjFrszJJZpYLnAhbdywdi5+YUF4s6
HBI0etW/akgvRmvBmHGdOO7mbNIVRAg0rvBw4/nRjfvvRPgeRdjm7K/2/9XtFRQSE661bNf2wu14
phgiE3IfvfKE/mrzqGg1zHpux6gZKj0rbLNnMc0VIJPpRLUiD8mBKmddVBXZTez+SXnxxb0Q81CT
Odt6MXLznY9q2XNXVYPCe0N/LATnqLWlSM6ydpLtNUrld+tqTHfXnd+UBS1TMvNB8zms1EJKIclm
mfUG3GORTjM7bIWtprVV99j+GGnBeScxlbaLVBJ+oWCsl+J6ywv6rdQekV8kiPbXasHr8CG/rouN
BooSgo/JWxBOyd90+jrshg/zUw13GyN2xL8IBWxhZHW0Zupn2COPeYEGsGnHpHpBRXy+MvED4pxt
i5OIsp+5zfB8J+s17wldqfCbl+mG4h43Q5+YWJY/ixTPtIQ/areOYhdUF1tivbvue4ZYaIiXPc0J
s7HUPMgtwv5pM+4pzczzC6zw6QkLJ78FbJODH1cXBY6NDZEfMHDa+NIIyrzjbEI+2pBGffprO6DQ
a/GZxOc99D4/uklAe6948IHLaTzpuTIOgdR7BTGCq3si8z5x1nBe3J7s8qd6NnamUUcOxipxKr1t
257sa62e3pS5Sxz59x8lI+kCv9g5aBK1dWku4yP3aESWAHROhZAKLf/w5yhtkoM0O6iTUAgtzGE1
fsaUQF/Mq313we8HPdG3HRGj+JDZC13y7lvYE7mzUX6jS+aK9Mle7NzDmr8mZRspZ2PRJFzEVFj8
KkmaGWu6kdxGe7dU4lWuG0ay9pwR2bxIfUX/nZilPsFOG7SyToQLX/9cIOwbVyXeK7HL/939Qlyo
uiU6sy1ejkUdY097hQKfHdJI64Y46SzKivkHqeYGs5ZY0LuibLeZzv7GwFx1hE11tDbbv6BCxrCv
0AXAm6YT88Ug6v02Pckf1zLU7bMOGoAZw5ryD2QzwId1yQa30ozt9guV/E2cjDV1MBEEsOs9KI5i
/JRSlzYK6xtm82ns5uDQUQ5FlXk2syIJemEXMnh3ww8WMJUIrmxSzlJfUATEy3H1A97dR9C1+Nt5
WIvz7ErS0HPdimKCddid6H2IgueGzfmLc4/Mb6HYj0iKUvgghnAy3Jhu1E90G7FMBXhOApRI2OKi
4j5mFp3iE9T8+uVN2mZVSbLhUyGZEKV80dM1kxY+Bj9ASTrFpcChqiRRfhdzjOIJxAJoDNHLMk0I
8fblpeKL7T2fvvgh6OjwbkIMu3oQ9isATJvFb7Z9de2TvSj15Imu8USHn4oJDJ7KwZAdleSQzpKz
YQDJLSHIZ2G4dtsgWBJ6lh1xnIkViYuT9umZvFdj3XfB+y5osqqnv9HkyBTF24fQzcLLNAv2vnn/
63zqO3PUzKSKDyDD+L4zY3RNMpfRRokAQvhBjPVQ54o2tNng8fhrrusAb82BIDjbbSE2njUdobrs
Ceim74CvPzB/gfSQt83/dUHBBuTZoPvPMW9vfKjNvsqKPCD/MLGdoYXRzn5wI2Z0kHAceG+26AlR
PcZC8s1q69oMaOno0YnO9ENFx7Teji03mrpZb6KTTQPbPgNMfgb8wLF+mES2DU0T7YZ2nxh9YCoV
0+r6Q1tTOrMx9k+5ktGBt1GjgZ4lgmVwGrc5bsEWogT0vH2RCJWkHnWDHboBkvDDZlDG7bIwUBGM
n1KCDmlciHbT/amuX3r7Hgk6c4f89g4dp6uCFbwSYqVyKZQ+ZtAH927QnVk7cPwPqJAkU17/9LhG
pXx4GL5Z51YZysqZyLGiPO24n2ajlmP+5lYwcoo9GPwwTmbZZRu/HwpYjRNkrKGs8A+dRudD498K
yB01LB9sw+2+1xazj0pSpHJMWLef0Gr5G0u77ZWcBMwB+M2uKMr6LtHIjNoM9h/H/zlrp5EHAO45
FJVyRzq1VSCJISzT8i7G1vs0paCdgL2ZgQQGZkOPDQI95wTKOFqolRCU/iKqz8ba/6RYIGe6iAiq
L56QLv07vcWObm5lriYIkxCpQGhArH6dQNKSajcHyUcGNWgnfpIDiDppmMz+Q843Z2fYuSMdsf9t
PVsFlGumM9LOxEZ37+gs0iwZhjefBJ6aUlf084Bgo4JBSsXntLjx5T4eY0f98sNl22hLqRnlQXfT
5UuDaSOeL3vXY7qKWhZSS4HIXXeWEkNj5bEZBOj0vjlq7HOiwtSpb6Wb4qOYeu9FB4/XwBtDchzW
ns83NvnHTWEoXx8NSr4ouXWUUf8wO7R5s+JJ8xhIXTkye9v+rY33PPtywXwLSd8Dvb069xi6Bygk
0+OjTU/HLprmMG4Zu9LLdjHgMHtZgcldy778osiRppUqIa83WQzhZCjQg2gD1R07ljJbLsdihceb
N3nTk+98NWP7cqIGYIlhezgNwhzDK7ech8Ak+mqBe01NFSWgG7cYs3S4nf4Phg9Un3Ip1R4nYRxc
q/dU6ECBv04pjWcHV0uWDyVdsQg6eZbVqgWsCFDqc5h2fLuuPGGBxWbRnFFsOV/tKKQTDwGffLxv
QUxH7pnH4SEJvr9GxcyZqSSr/QFFL5x16ZvPiTExIuZctb6WjKIBB7IwgBxBcz2bdwVolEcNBEC7
NYyAGkZX2j6qp3mFHTi/kHXDx1PE4YvCBWdSPQqdb+Wo0uVthwAtfYCB0ntTQgs7VMIC188hB1cg
62eEQZ9hSkP3MkuF8wm+dCbUoKIkkcE1fn9iJtJvJbMKEj91o/Uo62T36Agr2oXPp/1A4jx+6Sl6
QZFAHyyEvIPuhHHkGuU2IsI70T97q3YGUlRtJFluVGGsyS18MOqgRpw6O8bxhiJd0Nf57TlbsiZJ
onhl2vgVp5c2rYWsNghIdssoH83BB/lJYJJo+x9QZp3AHCuQHhziD3V4iauha17mgsMZFX4izgm6
ON7h5RDVGytytaw1omk4po+6azVUdCciwOm08w47iMFHpt1vKq2LX4U7mKQQSNpYFQ88xpj3vZnl
gSdVwhLXvYTQWl7/3LJsKXIe9qC4nsQpAj5a3imYpFw7vu2Q5WgBoJrH3e/v9WnE5juDtBXNXYz+
7RPzfJpm9BHqOsPCI3pWJM4EtFJY4Jz6cq0IZTwtWoPSDQfmUsi8ZYCKoN0airUp4WzxPdbZgafO
dEegQnMg7LycLnYB4sZR8e79I/t+JmKX9DRxfdDaMuPpXaGMVF4jk3CYUyjtNBzRsUYUkKaJUPNm
XafvjaRH2xVEPmG9pMn6YfmJHUWlwg/1W7eGiJl6FuCVu1F8DKsYSJmK7GiN2w07tzLNKI4O8yiP
GPEFLBGk3AQUA/74dyfpcugtXCweLK2trVeC7BkB/bQJxs5CjcdRbuPm+6q+ZGqITXNsFxOleY3A
uizaYLBQUsuGTMQki+EBr+06L9X4hOZ8udv7ILQtu/sjQe9pJ9aCYQXS9RhnjtQAlSWVexgDzTmo
+EMkRX8QEE3GTFHTBUxer1L7aGfrJsCmiP7pPz6zs/6nRNQc1m/O4s+MDaq9nJAb2pBXkDmVT6+I
TL70Gw86QbTOoGoHTxrjJedx0JgdPxmLgCzsxPM1VJsDFlTlhcHbB2lkLWJN2eKRWQ2isBYH4oJm
S2Mr33IsBBpd7rPdjr2HeO0/xMH/qi2xxElyNJCI5x6/hbBS2JEULvx9R3xZQA7/kaoOJ6A01Zh2
g7viKELYlmC399Z1ofwiqN4caZdnQdtYwVPei3FNErXEF/N5mlDP9tWjtyuWDBx5X2KX92GdVtPl
CpWja9HoLMhf/AQV8Whd9IxzxnZOCmmeiW9NG1gAt/yBsDvoMRKn9PrZtpeXbGawabuRhOiO5jM8
gGwk19kF/cMpTsrK23OcJxz/jhjpF7tvAISaYjJzBs1o2Q3BoQnV/Bgxp1HBUvZsaXL5okZynmbx
tjltwZXHai2HzAGHYDKUDYl3v49IAsNRgzzjjP5T8l6KLnVPGNa/dfKo9Tb8cqLMdPfZj3mcdUdq
HS9ipAunB9+5rYGQig/AhD3XrZZ3LNnHlAS7IwHTk87zmjrby3yUK2beAUZkxdDOc229A6gka5gb
zdqQB7MeVWHQWJk5oIZ/RLmEnI+y/2hQyj9Zspb0P6OS7Aa1huBRbHKalKt86fUgRFB78I4LPyHU
xIcBLP9dvoqPnB0C1e0SCJYUD+pEoKbybK/0CNPeu2ql75pmvVBxKv1d0IvULbIadiuBsNYyCP6r
SrJevD11DZjzgrpvoAun4XF09ZCXyHax3vn5BUFXzfMR40kHdqNtbzn902n8+fyYiuaFVfmypfqP
KJ9ZazEVCQt8PqElCtp9XcRpLlHUIGp2pUsvz+lnRqwADo2xim8XeaNy7MD9g8BXB+YkBonIJUa5
odIk4TB3pLpSyFFkvlljw2ksaATHrg4NbS5IGt3Umas5cXWDSKSB217nw7vj47QJ2kwzEODOpglo
CnqtRWSbFiPiz1Sn2qO9AZ4kQ1cdmcebOmHD9S03ZCxk85XKvneHalS0fCXBJU7gSdS9cb3V4MYl
FZuDWTrCaxNUnE7vY/KUqjaOcBIlLlvmBX4pQXO2+BCJwht5NFqRExRZaujQGxBL21Ykw/CsoWNI
FGsilhc6Pg7y7hQkxEOMbWEpiUvVSbU8i70Oo6lQf8IhxjIi4tkHm/lkVC/DbUWrseqQJjzjRMck
aeBjflUC7YMM0XQVDJiSRfdHt/vbyKPqrLzSQxlIeETAT2oWOD9Gfh2LFEms+7yt0XRHGqjtELTb
MIubD7y6W3E96MfkpU2HxTWBk5qFsUc7U+H2SYJu9i2Gliz4HhFzGCwjxxC/dlAFbBlPiZkHtuXe
7IHvftgjh8Q9K/TINSi40zfMhe0kDqCl6TTa0hL8WDPjUjE6cDJGqeOf0qTDxVrGykSUx7mVDz3R
cpCWH2YO6XhXfk+J4Ruuy7gaNAEKYwrEBDb1PrJyDnzB0YGRIAqnr6SqEbAkOBXsKSUN7RbZyDOI
rHxXNcYmvMjcZ05aZztPrkdutYXaXspDYvwwP9EFlstovuJM7VnC5hVQkWJZCzu7qVfaATDeBYYU
JK2ZNMCK+v4zgR8h0ZToq6PyaTzfqW8kF5xuWONBXnXR45XK/Dy6//FB/la2ngpgQIuYA5tKsqVv
qOl6Zg2hWT5lNU7A/Ii+PSBrpH6Rm5ICx7oLJ0SlDhTrVOaQYw11JvfGIjuiGkqim5r2CpWO4ye7
b7PCjQwiUvsYymowOlg2iWMpYUA+WPcOOvhzl+qM05U2jIH+Rz8Sk+7NIp77Am6l0QSIiwgsdgI3
vJJbNxXW59eykJFHYX1b6P3V2uzWWlBH21rTC9SoAgojZPixqH2iTHa9Pq8zzc0kG10xw1kSMXwa
a/t0rllPP6W4cP8ilUOiEocN2lDfC2VJgw84qoMOsZQSOjtRmqx0BKV6Nl8h2tXH9ROtRD9RC5me
NC4puAXFTh44jdh3+n/qciGh6d7KtK9aA/QPxRWOUmBQRkk9DPbKUkk2AxWyenBaRD9H9WsgJY8a
aPMkDCnZ8QgBjEklpdMeH1m1CHphpolyahD5x2LIVjmpR3FhPzT14SDvjApgYUfecB3ruk+VRMYS
vfIKNyd305w2M6/t3//rv17tWGrnOL8+JNVeFtPwSNyKDXw5VDZGwEb6wqP3umG7BqQFr8UThcAu
shpvFS6hYStZq0LuqkZ+zBr9DLavhIX+kq1tiG5zsSCgfZNcvf94RMqZdTp5XKYem+nkCv57nnje
/i+2zueIXXODmkJ92l/MI1iLXkTNnKp8XruED6C+F5Zm9IBU+Di6gmgY7BfoT7Nqndz8qKoWpyEE
H7aqiyaox0lucs1Pb9TSmCN4oPzYgIAXdFc4Os6Y1jN3JD2ZjNacHcH93YqMMEAo6QAnVJSmg0Sm
aaK+9002Jc6fgW9kB8kVDSx8SKifY8lD+gEqQdIzwydtVSYM077cSTp5PoRK8cREmjMbGiw+Ssbp
jHveQnoS0MKQexPrcu40F0ZVjaNtot7jTUyQBk6OSYUJybTlqZngU99uqALuZ2PLQ/iSPRszFB2a
7SJ6lQfAs7sf4Ml3CmMfLMNkkNuR12LoE2DP7jdSdplZ/98KwDSjc0xkMHA8Wth7j8yjMKitMZ35
FAO2fkTn7ABpd9DZAfF76Et9XDqI7Qi2zLxDmE6rmtm8lxVGHffrytvOlxXNqyjxZ5FZ0UfDC1BK
XODH5J+SgoX7qLWUV3D5mqGn23ZPrIiX12FTt+5jnERch1X7YYzmCs/Ih3aXHWKDhYOh6Ww02pgm
pC/eUlM4YTidY04X/kVuU+Uxn+44rzEw2Lj6c2U3Q+S+qU1Y0P0X5AgITxsk7iJWtDJ7VqqCrg7c
W/cadEiejCoQoME9sm3Z1oTxNu8tW92Anx4zcVn/hbsdaI7+sDRq1nAWQ7mMrsDiwKRSHALBW3dG
jDE0+jWCGbV1aM27UWf2jIkEXYiLbrfBCTPi96cewZ+7V28W+O5uZN0CT21YwcR0c+vuSh/olFEL
jka6x9vtLS/alxKpm5XfE7+yVH1BoqkO75Q/KSbU/4j5aqIpNIv++qun9wYv8yYsBrjdqHDE+ORw
c6dQHJJHX7B3vWGiFlGEOBrLT3ANom5nnnNxDLIRbVo+AwFFIou3M9XJU47Tz288iMDKuUIS7l8D
VrE/SQgb7/+UCZB30GP31HRtECSrWemNU5LKLLxCeUaaeR/4MtYuycyba9l7O1QCA93WvWHeyMkA
pkywQMHW/0zyr8uBreOJ6Mp1/PGZ/Chj4JLhBFVHPHD4Fs4gOyFxqZcgq+12DZh305W4DNKH+FQ8
V4L8esz2X1ownVi3AS755iQls/djl0Q+Q3nqqfdS6ANZTa1mxmijgUchV/H7sTDuzFygtKiy0tRU
oW+u8JP5CPDn5Sd6ErlVeaafgs0pQSlh8kj+80L9yYGAYGpGDXo0bjBMFiyP8oHSnjPoVt1VcdTk
138JaElXu8r4/sHIpKgQYlfUkxbHb1mgGYDPp4nQ7LqIqyZIjsw9PYpKKx9Aq4Kupbj3AHlLr9RI
9tghOHMO1S2e6Z/PvyZg7zItx1HgaB2n9TgztP2QGq8SCaEgaG350/Z48gYsHcLLtuHbAM0JnrjO
apPPMq0m/LosO9oFhAEECdsMBYW2D9Rfoed+CpCQwF7FYgL2kDBq6ynB5+Hrj/LIuHuakI3YyI5V
E4e5NfH0CtnAYXqQxfvjM3qrp+sOz9+H7Qk3piZ69CkXGyNWvspoOdjnv+lVR4a8LJShGkJzY6HK
+IA3HK48dPf1G7d33BGhu4RMtPA7lhvkV9xgYGo5HB/ZKP3vU7r4/iq6Gqg3VBDicwH1aUy0u/tH
oq3q1EeeGxa1iGHv+4O7NJkZVmhqGYY1DhdDQ7SUJdRyV9kwaU2nTRZM40W8LA6LGyOTcnX84o4X
SzJIV1s7nH1oHYlvhYP+AYtsCp0H7E7ZK0ylpn1572X6iS1VVqTLZJENV5O4A2wW5KoEASY3iiEA
mZ1AHGQYCb1/KWaT2ADMgQXhsYAMuhvG+IH7Oak4i2/5PPTdZVegTNVTlVY2nWXUs8inIL1HYUSo
dIMDSiaIhuqxWnDzAlejxA41tqud7D0gE8IZe24fuoTU4ZNpBGtnroHyZISh5rY55rubZOoh9aEv
VS64N5D8C2wGCS0AJ/0YL2WBWXNPqXEKDMyb0G0oiqecQq1i7Nu+IBG9CKDIFC1e0MuLUjPnZcHk
sgmyv3Wao0o0/IV9eyzglMWAZveIL9Q78T88N/Sj4hrIWaXkDdFeUepPnNkFDqW2zqrd8Ol+ZbHH
26ix9cORpnI9rZ8TEGzBw6Cf6aCuxp/8VnrsplUijf8WVFYnd0eZar9Iw0HhgRAKlnmxRAKy5MGL
wvz4abvUiUeXqyNHxJIwr1spBIKIjSk0oRQt3OQm6VeisG0Y4HtsNobir+A8cP16mnloRBr8vnCh
oB4K23zd3TyjcaKBqQAxad3LcCrMsRNQ/9wj++CEFK4fy38XqwpD1LE1BDRd8wjXBzRbJdcUj8u/
uA39s+G3eHeIsB8z5bfsqWUgo65Bo17qCwiuqW8j6i3CwlqkbHzGKH7CyFBL2dueX/HsbgMkBMCe
VacMb1C387jPoK83EvLkGKEPt8B4rDHcluWmHIdxKE1Nr2Z41/vwNb0MCDHZr4fTauo5caVlHf21
aWuPpGfj10RT/eRQeK4HiTDGb/1GcapTJeNFzeauVJqTIQ8wph9h0Qi0+uktUm+9qlwmF74KGRNP
H0YN3j2s7G+ljBjsQ9++vnYifrm6Ch0dTMI62vhJggw0XFFM6ybz5yHhw8VPcrQtEIA1rbgjMBpX
KlvWOzmebblS6NZzoJJvHUfh+u3tvsBUy4KhHk1M9hfavBVD6AXoiChJUWQG6ymY7izjLpJFYLKM
9HxQ3sJfQCYLFl7S+VlJXFPuDTt5T9PcBSPMjNCLlkbcc3DAVMvGWzMQQEQW6XS4U5ERsa3YbJLK
OoFS6liLl+FfInl3hvG+1ruByZZn77bsmE/9FmvXZHmtplMJFpZz0Czx1WCkB6R/HIhaOdaPicB8
iuLuLDs8DMBMtzwi2oCE4Wn82dUR7uHJVAO/LscVEBB13gpW9C6EtdTLuGV3JBZclVCf+GJ2bl5d
p+6Vkx6ffI4KA2ASSNA6OBOI/njroe4ezGdOmdfxbteB0wRTrlUpxPbDhBefxTRHnCqfvXEipPHM
KnF62+CpW5KPt/ZAoNsYLdF/GtLfxZFODV9vG9Xu8BoMI7/m7yWxNGwKk9tftmeKEh91lynyYNVz
+fyKiGxxGjyz8i63MagQKyPZHKp+1gyjz92sLRzMmm65FNEbzS1gAg/pa0zEG3a3gb0feGqWZqLG
8Crvy1AqpL99dcwP+UClwxJlDiumH1RHkLi8guQZvqnnOySQSZjoeQ819p2B3tfC+ivcBSAL9t+e
t7ETExZXFsqji9ho/GpgHwzkHc1vHMQeiuQ/WDsaGxj5Rmw5crMFqENjDpCDoWIaGDxxeIBqnSdk
Bg88STCW7R9K/fJGrICRXqE/mx0B14GOvDrQOXBVXCUM0tjxkNncE26EYoCTEfmCPZYvMmO+x6WF
ZnxONAK2qnW+dLHDFsPOCsumbRTZAW7KQk2RHKiXNpa/Wj2UjBKi6RcBCW49/RrlnBTnszsJ3AK7
p4B1LOoJf4pRkdbsplSpzl3KCfZP2g/QJPp2zhtVsZLC+WYfKab3/SU+mwBInX7kZxKMOXB8OUyE
x3gjak5bTfai3yOra2Bn1iRD6pc8qsTkGnU0lSZHxpskKNXATd1kZL7LMQbzJqEX8cHAMOqZH5oJ
KmKT9qw7T7ymN/v5SqlKnexmoB1Ewr1arId6jPtzy15Ryx9Pp+UJXgh4/7x8aAraW3DuNj9oxx7i
tWf3VQrYfdwD6knbD5CNd0To+jGydn2vF0bU4+kqL6RgbsPiN7jZVA+RFzC/PtMajr7Oa3b71Ykz
AIERSA8HajpkP1pif4By3Xh7Ceh+dH5nAORmIkfv7eJHjNGFphFaNwMbAcP11ZIqsCH5qOixZNe2
vbJGG5vXf+rINa10J5oEZU2qRXFd83S7e4J+Iq32QFqLTg1KuuHmt0x3Arjvpq0uWBUUHog9aYwZ
UIcJmAS9DyxhTthfYIsJVCOP77NbmcRYZg/hLa+UaLRB+r/jbA1LUjgwfhIsRJlKfZwnJ8mRxLbv
I8B7fIeq4Cq7dA9ygQvwo/GyLkOgzSHsXTqjDdFHTPOFe4tFiawQvi8Lmy323pk9zo2LySKdhPcR
BtyeoNzf90SlsU1txOYytA5uL753uVhUBwZ+9LEqH1FWVTuAbLcAIoNEp/RE37ISf56fG1+oQrnf
3jn5ZkwwBx4fxRkAKwwnHqzGKsXM+79aBrW5HFI/G6mSU5STHaRaQyjXC+lhCLW2KIon4J6MOJf+
EbmIRxCJmK6lPTYVAGFlLzFRTYCMD5rZNOVA0RvI+PPvlJvRpTCwG0bZhyBc7SIXE+FVLzkJvsoz
INfn5tGGcoA5JRGCOXsgukDjG+TW6hUGS1Z8BX1IoLZCiWtFBhSUMemIBH7IzoyrUXuAHZKB7Djm
43aUbTzMEeC5oWr8ORAScqZfpT8+tvfrejXR2k0sgpl590Yr5qBqT4JzzFoA+aQsqQvAa2pmRbjC
Tr6LXrvxt9ix00792wzNJieNS5jKw6K+SGFQKOOOVTBFi8SXMqRMxxRGdNrL3FYHT2N3BQkEJpeN
WpD16/9kUFRlbTFaaIsHTFlzGEhH7sIiuv3wEgGUQJQ2QVAAK3JEt1Vf4lak7dTkOSoyyClKIoNl
h4kKhSIUWPt849pyv6TMM26NXwJ9LfIr1BBKefhS5nRGQ3QjrqQzcldUE0SYQnDmLKlwwoXmxFxG
MEyW5v0vtJxGTyAS0XI5tapT0ZPLdYtxCODGfCuZbHMHC4QDPuz/eSbWDImMT1B9Lk5dAhCdBZ2V
H6+VhErfAmPV+U+ywS8Xrcd/vM5ma+CQKBOf5k9dxwI9/uoy3APyrU085ERnImTygQ3Msd6wG9r0
DSLU2sCMgcphL2PbZAUeVw7d+TAR/UFxa/Zthd3ib837Qx625dEqZRsSH2eKysN88L8h0mvXDZJ6
luVyXQYEBr2SVlj6jW/HGHGIRCR7GqSckzROJmnir6MUj7imxBjkGwB97l+c9aN7qvthfW1PID7j
k48weDLJOfQ1EkGJEgxwNOSTduFoprqZos46AzoG5lfSx+nOXkCKherp1UUE8Uy1q67EYTuYn2VO
w0cmEuZ1qq0oVST7DLa+CzOp0euRvfKzh3L1oCnDOTNNUxtA2ELS+QamOc+wT54MfK6c+OQddn1b
GrS+clsmL9ZLR2P/HkSAeP/enu0HEVZxApl3bIIR6nszBkZPPWDvoqErxf+Mcw6SydOXe+Ea3C1Z
KbYxQLMOTSiKGvjeM3bRcvUgVMVoPW6NPnZcYg4FYLdmvcz1gHC0yb/4VIm+H8nZeC+JPJ/JlBWh
VqtUrxjJ+1TN1V6C4Su9hRTxwhq1Ssjh2XyzCLF//VNTx+WRQ2UoI6W7D8LiaF0rLcyaznlpHP8N
Nnw4icd1cX/AfSEU5TwTb+cfmzYh8IQgAm85WTi9r9i7vfSRRJ5feQIg35YXEM5G4R4QWLcPiw0B
bnGWQgF91ojxs99Vr0I8oGjrBk6Wdotpggc0Tuilu96WFaW5G7QrnZwqsZPTmYjEzK/croAp8jLw
M4YyUH8L8yvgKjZD9qRzl7HWcGw0RHQEJ7aTNHhUPDooN9QfzYijPk20tDVSuhJq87z6RaaEdwNt
oD1cZ0d/lXmhvvbnikqgivCTZDh7yqV/8KL/gN/WkqF+p3cBShoj4ZOKGQWAJg9c+TEsHNFvZJFu
mzMECRo2V9Vjpclr8Jxo8i19A2/XpHjWEQ2zFpvNkoIg5r/CWs9UPeRLBYTWtN5qEgTw/ZtLo78o
vSnVwiHwth4Y2MbC0wxAHRRyOLSgLo8coQH+ng0qxEZxLQTOixsVUBG6FE/87W9Nwmw1o9n6ui53
GjlQfw4C3xDEy4diVso/1uvrK0lexh6drGCQeG6RO6QMwdK+YD6QnXxevR+OV5uX2oZU7NQxNJvJ
TlXY6pFB1M2Ck/cPKefBlrtE4LMrGaILEaQUEuj1jpfrqw2wMjw9fB6D4HDN+MEDBr87j2N11n7u
EEoykdniAyiPRHDtoGCNrJyLK0w5LT+EOoEocnO14Z6QsriEWUOwXLKi2vHw8heGSqbY0NGoNBZo
jTUB4oVtGtatLM3UFp6uoiDPfZrd5jOORvjXWYWoK7qsiuDcavlMqFHoT9U7u9HxuP9EwZESoe1c
U16Ri8y49W8JU+K0RiFIxmxz6NSpSifjbUfVtJeXjZ9TOvRNGTgqs5r78rTKqn3inhbkUNb8PhI6
p3c4NBjJt+2inFmXstR2x+RPUPAb/th8w1oMSKiZ5VRfedB4OjXvOnDIPezpnQxms6HrdHmaDCsy
gPUFnt1fxiR8Yv3xVh7wFI8dy6ZGmFLblb41RhcFcwTclS1G1VBMdw22n9MpQjbAUfIe4X1ufnzg
mh7RpaWbydIpkgj7wEuMmK43siEXpkRZ25XQeD2VZcBuCMbCcUT9OfC4egKY92OXpbyzhdzVA5Jf
7ZsXqRVBiB3W9ac2w8YVlauctR6snu5jiDTBSAakEM4M3U1lsSWzDVLuFCBevxa91Tcmca/PoM2Y
4mZSq3X7U0hMXj3RFJTzqD7mWkLNh2lPxHS1emDRl6ZaxMeJ/CQ7NRzp8oxti0fS5vU8TP2WsRe2
ClIPuKL7AZMbPCc9gR9NUIQY8MS1gqzyecUldRbWdZdZNIf+BPzO/CfH9TZEZmcMDrRyutlv1OsD
cJHodZVlUzLhVyOqRFXerbW+yt6lKCW44syDODcRoAHDTu2pYjeIW7rLkYtEd89bol4ywMi6uKZQ
sQo0BTw/X+cmpk5+ad/hOkbVntU0uBnuw5wab0BidcpqX6F2XHLsPzMztKPQpsIEDUHJWgbvlxrK
EVLCRM/evz6Xz2ZCVM5LxzwR6rLQSkVJSZgw6pkLcvjRIxvuzn2Vtmc14wKN5Qr3+jS3v10RGtSy
ZIAdxQGbihC2fdiHPLY1+lqBXaQthhtVfeQ/LIlFogCkmTEEXll/IUoWioGdMaQJ2z88rJy9eccP
i/fh9aGUIAnG8XYwAd6otxIWFrntu1iK1FDV8RhpgCHKucoUxPR42dAmp2woGDrjREsrSYF3jSAd
+DAlbOF9QEXxS6cyVFoFvI7bjwk2/qJkF9BLKPhBRxTbT5NTcaAt+ps3Y3z6gqBkgGsMKePIuAI/
ff1xALEhCavaUtLhBy8bKx/n8A5cO4hfDNzc2EMG7ZP2EwnKHmTHHXUV+DIW4N0hQ6vGzERRse0B
zg1IsbX23ESna/6BsFsaLNKOyMiHpiaajBbRKcPmDvcfXLnhzhWQe3uZg3Nk/78nafxeqqupNFLz
u2JS5TMUZpaiim39ua31UZZIzbGiX1dnRcE6L5t0FMvPooMBVgzpsBz32KGwzfl1bv4GNNIsUyJc
z13rrL3Be7Ul0qIEfLOFc44ztbAYyg/QKjixRPzBShzlFz/30968ZtJUnkoxaGTaJnhb4XxwmIpU
0qLG5OMi3zOq24CL/L/qF1I0R6+igcOJDrqHZbdnfUrYJKxzHYX/IcZJPqhYSThWlzHNmKiYEaHS
DWFvWD2xewnT648+328goIy+oRU7iVAe9JWYx/QY6cxMCLcvuNRq+p1FqeawWO+uOSIZ8dbbxTjZ
hYXG8IgFSQ4eQm44Z3bKC19t3LhDyIDY/OEOErXJiaeU2dsuiwgU8Vo061Zdkie/Xy01gVdDnJ2F
Mu/Rr+jHLfthTbHePGVGR/lkrHlzJLqX6txRa/JX+b4wmSElrNDkJGoeMQddyB351oN7lS9shIe2
pTrvpeGcmNwfCTyFw7uRyCql1qcLo6udTeL56jXIF60h7qElH8hdMjNOnmFx7iyHeni72rBGRCJn
zGmo2mSaCzo2zNs1FbjJlq4Ja7y3XzER6HTTFcQa+oPMGKnFgMzsp5KQlhUNXq2S/G/t31SxIUJz
o3tjoNaGSMPQVAadTSyeXCF6aju1XICwePWuxu+dDG5TuOW4RxqGyzP7+LsNlvI7AFVzGpWLXM6O
Ftrr2OpUPups3gf9NpmdJNPgC4iU6xmJXl3OaOE+1JDA7aMTVYt819k4SYYoIGBkVootsT4EuwFN
/0p+ALtkKryH908jZ6ASoBMtHp3JMsZ4QJaEe7zjCMS5QksJv/f6idsf6rABIsLkOTdSUX3ATm3n
RhR4XU/0Xg0J/xOlrlY6+mJffIKr3UAovP0lqUeRLmkHCBD1ocVBbWP8bxAllDQDCchnRi8rmX5M
EQEVufAkqPhm+CjIQzoufIaGg49BaqHYcUHeE/IFDjDOpYIWwTWar15kEI4/cevLKOgjkrl2KZlS
xrZTLqq9dG8CIHaWaUTzBQd830MvHdMJmEFXF9KycsfW78yrR3tKxKMzZSR/6vHYKL+8T7ct6aw8
NunsXK+8yKJ6Qt2ICVdKnPci7c+VBLOaXTxyKmr+9VaEA1AUfMoxSr30zMD8zlu+0/cxLN0rjtxH
T704SLK5NeaDbnmw+LocaJexP/bG8iw/Gh8p7MRYpD6698NND+RCMj971uuUDeGENCHXru4lz/gh
aW1lM9/GVGE6w672F3dsEDZtOJhR2V/sjI2G4xh2VcG+cAm0T3t6CKssZRH83PC9nQKlQuafVIDa
AqFay59YAb2P6CjaL/tzLPh1fFpz8KBbOo450i7VIogKDu0G8AS8LYWhy7NZF5D8FP2CV4WM7nTG
xH0yGZvbSgPuUFbq5Vl0THm9mgbNgsQjSro7u0/Q4SAUiYPayLHFHTICyq9EfxLuS22r6bcZBWDg
JxZqdWHjBfbyrJgQ50IBmwxi+T4LDz+wUlz/LNZPNHuSfdu0vvHRpF8w55gr3vUEYILNBcYJj8Hi
8MxWQiAw6JXhlWsTkC6zMWusur8eBGZ6ToD0wqgVh2b2HiedVG1Ijrt4GOu4Kvx2RhVsW5L/9XKO
fBpRuoSXvSDhy/VNPcE9jsBr753pTw2+lhST5i9ujWFp6V7FbB3j+xRprVZ8Cqwvj0RGfHFOrXpo
WD7qLJ8Zp12V4FU2ghW5J3qkCPRoMw5e1GTCVks2jSLir0luTNwtkaZJ5gJKowS1hxiCiqMoZ0yC
Z5K82Qu18XGrpjxD8C9MMVIlbqQCr5b1wrwVxXv0VCSkQw5am9QxukH4fbBzEx9XOZG5iU8fSzdS
8af1xEe68EIjx9fFZExXapMCT0R2XcYB7fNeUdpedKKEhXlfIxMiFtTxGyIm79LdDrVcz+UHSbZI
hsyVe/Qj9QNn9907P2OJPe0wqZAaUAMg+fxxqaB8SlMzavuC0Va+tRsRrptTI1lyY9lRgwmQsLJu
ZQeSl9fdcX64ySIDpJbfJPryXJYLaijZZw36d8W1Z1ieJZM3XIcjiw2cX02ye38ku7Jgc8ZIPwkb
Cxt1h8+dwu+dgxIJfl3YLvZZuRCzpg8FIvbxUwaSqQf4/IIxIcbvQnRzq/TXW0w9MGb2BMbKudxV
88M735daln6eKI4U78qvbLRN1f9oDKZ5da0EEnyYObodQ8LjaJW9Teq9HvjydKm43ykNWK3+Savd
4T8O11xaA9+w2e293MviA17f8R1O8l3w/p1lq14cgD+kPon75UOr3P7o0pvrbSdpTI5qeWdieMEt
T0OrWDN4bCdvJl/7erPnfIUD1ACxazS/OtBStMzAchvtj3bnfqrgZxy86bhLrzE4533DBfpGJfXo
qM5A+oSOOHRtbZiWETHecxKOMofhkJHD/agL0NvABF2lEjcuZ5NvHF+nYSc+3SM+iebFx+W2ky2D
+dNJaRLt9I2rKfGYfQkw5Gf1JML4/U1Tnw+GXn9UMPnpSdEjK5owOlNUTpbVqbK8rozoG5em7PWn
p1Ui8py6iV4wgnFMCD0MgqGvV/8coR/FnD16ZAXxd2YhaZY4RxtPm1dAaoULBVerb3V38G+VJ5TQ
OM0MoemiGykaUjl/4VzBvjK5dlm5OeMY4S7TBPRNKO8Zz4oNw61MTwD4Nb5JtT/pzqC489H2ZoFw
+WMGrulaaCwN8UY/G4dIYHJbea5l5G3NePkkkm/osB7hwMMCr5EWLvA4al3SEFEum6jNKP2xxpxq
mruVFY/pGIuasZYzOGPOIw0q8HoWBG0uGt40rysW+NhizK3rCvRAGqAj5ebEO+HlObHlxrSSTZsL
M0fgK0iyXw/wkq5TOL5+sRNQqVwH8alUePBRLZUHsuWl1K1gAGlvY3Qg11ijb0/iKVo0+3PlJdUE
fm5Oy2jv4sWQgEB+mP1x1bEJlxVUf5cOFbEfiCAnJaKhs6ZhsL2/CnRgyutHFVxrb+LraQno/7gz
JMsFp4dOIAv64zdeBl18IBAivA59ichdDazKz1W2GHsEWQjofd48/NdgO+QKi89/9Y0qKFGO9e9l
ntf/BMUr1SHdCDOQxh8j/pfOCk80rZGIaJO/bZ2jmN1I/A5iTuYdAB3I21/g26A28RywkQqiX3KV
aZuYeGf9NwFJTbcM7NXcLDbV3aUwBGqsIQwk/z/tX4xMYNS6H0P6QqoC0uTdDGIJ27neFZg+FoQi
qvg/ieT+Sktr8mWZVOK4mdOC77tEqkg6p55yvunNehiIGaZv5n3a5vMbreIWV6TjsTb7q9xKIcQA
gWFYox8kIzNrAnIkxWsi5S/ek/SQeG+g/CMULdiUa/YeHPzhJBf7QYqhiboYq7Xvr/580ZXVHywn
HutNsOFXAZ4Nx/4LuaekAdafJ/KzM+IoA6GaQ/3ydoKfbxXZHU3+9hnixagdlMEsgjF2Ak5coFbS
MMHe3m2kDgn/nx8CpfC0cBxBqOtJWElpFGWfuitZfKpsOkVV6jCNqI6LG/Mz1MkpEEmGCJayh3+d
3DSJcBVwJWM4CnPHI+h2XItbBpW73uLR7maCsoCwVo7XyxdkQIe2awJFxkdRErg3Ei5hWkPuXKNE
HotnIQDrph7vj2m/wotbfod/Vy0ffesbGqgAj2uf9a/GTOWBoQTP4G1/HehyXGeBuY8Ui8ElSTcY
WcVRxPcSXmngbuZ2mIfa4BD5NpRH8UgBogtURYRXcGxztk7I3yGQj7gND05oDIkQtibx5d2LJ74k
gnaD1VNDDTQRGRaea7docXy42SW5elF5XHhgAMMHkoGjuJxBDlLNCRrrKZgUBNOa74QXbBZuJaXI
SY7i9tqAuX0X513ltNc1tf0gxApxJfHGiqtXqcWB2T9NWNB+QggAM9WYDGgJN3lr5ruCPCwVOQbZ
7y0NL/HxtRuDmyExaOzEYfI89uPS0yCC18n7zrGEnkq9mk5BxmCSCRSCO11uHa4uEeAHhB2JeMmO
mNkEhlfEnIfVZBAZ0y9D95L/74j9CQviXu0LmSQm1FNViYcBzsm8K7TKQdBqVtskOiyjmKGfkJuP
FYuhe0t0fcyuRM4dFn8rnd1TfhN4ZO5pHlPCzb+EemEjvgR6iOiiEkJZgSLbM1rqJ42X4V5H+s4/
ytb3Pq3jxA/RacdBL5w1E3U8W21imhtv47nAnR0SIMhD/qxzX1aqVacopeEQrYXyLzFh9+TXnt6t
oA2ea/byV0PL04eE6ADKI8L+/I+bHcJmyq0RQ9iW6D2UNC3tSe4yjQLX28PFAJIl8ArY8TBSOsaS
9DhyZL7dfZLgGBDkMVnOL9ZQCxc993sBBVzPWqKcZPgEYSk73ATiRqdknA3da6/XZBc+f5h6mHVJ
XCstGqzxn1d6zumQ83Q/elvF/uDCdsrpbukfWjQ+lH+EjoZ2rOZsanW7/Q8KliONxskLIqeAFnr6
xxXqafUhb4hHImAfCVQ28qyLenob6s0VitraAqqENOCQk3Pv/JxaUZkI+tH/BPcXrldXHP96LoTQ
vsY3p/JyTeYHD4BFWNQ3EWtkoXSos/FRjL6KRN4Jqv5BfScRZurV4PKeZE+K7CytDk5XTDlrkKjY
FkRSDYuJ1dKQMocoARw3vog8RBTMtMYn23+HBchrA8vTtjXorUzPlFTDihYxZmuya98UNd8ciCDj
5ymJRvoapT/AoIn/OKGo67yVHA4SSda/4AewLvPy3Za4Pd1Fl0A2GYQuiINEX6VSeLaGvHeo5rMG
SJ2Mt9Y/9c+24Or+HfKYKtqllE/peHmGkXSuGsmNro1DIMfOi6xZ4E1IZgSidEmeRCEnTnt4gBex
cqzdSCvlouEP+FCLpxSmI4MkRruq9o6OANzbM2HK34JRH9LEPftWpiojhdV0NyfShPDcZUKbNXHn
k288MfUmNhIJOYsXf4KTyIVniPaNyyG2YSiW5fuwBK+UJ/tyNol80eK5IpvR89Boj0a0GKGKQf14
ychEMdDUSbw6nTueogC8bqd6dboybuGe/KU12OvF/sbl+y2+Ws8oQOZ5UeVHmQZrnbAy1WDGlfCK
1I+3z3FVOrXYSlNlWPWvaTGeQCEbc9O0cU2t+eoGaM5ZccEPx5f3Dh1N2UHyAb9DJNw0H7N80Krz
Vy/3T/HPyZkyeBUk9jgBQYFp5Bh1l/aiDmOTFLHdx1nY9VJ55sHLCWehmddglr1Tr1We6ir8603w
rhm7xCZmNSd0GIZepC/5OHGqJUqwQwy0w4+jy+Z2Z4J1vaJZIKkcaGdC2yL79PPHtNJ7IaU3BPo3
NHR+qRB3O93kHeQh28AMq1w3rXgHAVaGwfR87VEE73tuMPpvqUxlvgYAz7foXI1R+op+YvC3DzDC
/yKS7/6hQ6LALXqdCJJhHAwvdlDOEddnKEuXYE0xFLORGFUq+qIP7v7BSCyWXNVGGCiV+kPGr5KZ
Ysy1INBoXX9Gz8qaMoiR4aGpxUn9elhMv8nhQu0DQY6hFRbYmknyjGGIijOUO0NrtIJteO/XUrZ7
cFkykF+GpbdBKDNajcQNOIg9yma1hFyFOBC0+gJ5odFrtRlW3iMh/E9bUSHhcnEi5/n0nci1HzBW
Yyp7Hse0dow2GyjHrimF5CbLxYtsc9UGtpPHnRDdXn9zRciOqaPdLK7UESCe17OIh4/YI3dTUtZ+
NcCnntuCNHwhPoWTT88MlTOzKn3If7XhP1E5OpgkOeubQZ7n5/rBOqvxkSgIUr2rGu+BnmRbO0Fc
tgOtJDSN5trUWBuMsXB187RJEyYQfIMpoY0MhQbXU7y1dReM+LIdnA3Xr0Kmt7J2rXINkieO8H+2
t4qWVMrx5xbKZ8ZClvEUO3UFyXPBbjwEOgcmrXax72PiUcY8CHTHZTGCV/BjPS8Z7YYB4M9QJgwS
xKAetDN3RGI22X5iwpgTEU2dPXFw1MRPHg2CTy8ANyJ+6C3NMUIvSrdkmcY7MeRbnAmnEu46aiDN
lBkdnBV531wN1es8VZXdU6phwxJn2lKB3udVtmY/qsmxjizcnorVcZvXrGIQFuRvzAKgyY1JBm4/
/zBCzAa1C7UDHiqDzaEyZEbI4ExjFU4cLJjGLQ7Ly8klOu9R3NBavA/UVE7z9syoosafTSbs9/8m
QIChsGocJ10PlMU2Tbl0pZmxesYLBh94cI9VpEjfsG3vQtp/fAw8e1ehjoAAKEKtSJMlfr8cVKRL
WODC4DGE0IS1E6xPltFGupoVNPpM6TobP1k7bwe23s9sF4cPtGoARZSf9OKQAtp06WoU+sGxNTWe
DoNsYmOYvaMgA7sVXudg2gcRrskH6J7ogqrJodT9CmMuWi+f1/qIp4MZOip8Fzu/6mcp2UPhu0UO
0IhX/jN+SeOD4fSrXveh8lELSwlTJZUcYKb6WVIs8cd8DWMRi3bnZa9U/4vU8DdRgMbOVy8YPn+c
tLcJYgdPlVM3mYDgc/R/8MQplDnQNWhezSl5HkqnJndp6QBsfsIJICG8IheTICFnzgUOvFMSNb0e
OhkLUALH7pyaY8oPoKMvZ7ANP0GsIRIvcRkO/e+kvQZwlqmmZYYmRlOQ7agPKXsyz8Tq5RUWovi0
jRfKBoceymdWSxBiV/FuWYEXjqTGZWUXg964pYBDlmnn9VV9Zi1Air/9oN3dtHw2b3oV9wKpN/qd
s/92qVPybM6wfcVAn/ifNmwAN38jSWEYslf7h4305VlEyR2tA6eZT2aTYxyfKck1ZO2CiHf23ANn
F9lXPrmSQTEuOBGQxKVO1DxX/CnJb+vcqbyUH9Fy5xZOgKEwPYb3PdFKZGsZerkcYYTB7TbxItlS
L64NcF8zsT4rwbgu/SgYY64tgXLt7KFdMR8Nt4CA0VZ9Nqjj3u4EgVSd3gP/ikcZUmd/ZD1dZg86
EWECpV3kkxXyAmfMeDPhbNIJF4+q/jBp7lDXc+BdH938OyFfLf9Q4Cr7y3Hm0rsVSK9CG76JZGGg
l/d3Hqk4Mrijn5zjnpgj+QEgc1REOWv2W+MWvTXus8e8URDntx8mkC8w5u8rMt0yaU8q9NoqAIi0
cTmInHvY0aP2Q31voKee/PhNO8rT7tUQ1/ZA38tSn3nAXBPswE9eJr1Ou9rI8Ksos6CGqThPxo5V
TBUdwBOvz2WSL/lBj9LtM6l+SBa3wDPvvVHXfCzjd4Ck8cn+jQXl5Ggg6MVXcsS5HTBx7JcTiB/t
T77YN5Fv7kTvV01EpJJmwnZOXu8nB3uYn4iR8+8PkYsPCHIfMXYm3nAh+G2UP1VUXgqJLxFq2j0t
ZGk/36r89H9o9kQK2K6yei+59JItwrTM7Jdg07ZVZo19owPHDq4umL76OToxmLs5rqvr1fEyN6cl
8yxbw2oLRr9xNCMngeM9hhwcK1/B9PWxZniT4mPKjyQURYCbMVtGEL90lDx0a9dC0TWgEyvItbuC
WXBaIJBso3iUDCA8erR9ssbrwLTux/onitEG7HsB5g0ZHhHDUmnwHUXLawtpANS+n4HjS//bBbG/
7G8MepefphRVdsT+mMm7Qdn66xQlkACE/HFRzY+2yDDPNkfr/gvAD3pXFpUE0tdRkbJ05Xx+wqiC
YQYMBQsxR7Y6quAkHu8c8J8fpJAhVoR3Y4o4Mljvp2oep3WgOc9ai9XRwgW/0lynsCWxc40L70wL
dLfHdxZcccl6sGWgadUmR0SjbDzNOtgQIxfoFdYE311pXpDrqU9mMTfM+w/8h8XmPdIw1IKTzxXO
SjN3kuW3YE8PunCFCRwIm/GLk8DLrRyiMAwqFQUweaEV6AcUzwR7jDLQvvlzGtxcvcq1PydCBa/T
Bkb6eDaYEhEpNNIBa78O5f3TcRVsZp4BN2mlfib2o2IlwEOUbhMnCaf7YVkvcxYsRzoLusjrPf3G
jTfa0eP3unioEZtyb2d01gL0VXAmlWTH2fYyu60gbIfaDj5UIfE4Ka122Avc8DQ8XEdbVdT5XKa0
XSCncD7AZs8uvQVjcbd4P/Uanel20ACiGmpeIkiHIchAREkzY36TjrrPA61xWuca7n/8IqUypxc1
P4u+Bu1SfdAquos7VOwRnUpnxSRUGn8wVSz0F6wQLfDm/h9C/K3gIB85oiUTxXf5gwCTQVRP3bOs
JsNSHlgKe/7hj9eGgwlPDO6njaFV5nre2sm5myPLUBdEb3BRpleeTFHAudjGne99AbYaATZrAUXV
+y2f1L0+k4sDxftZFb3MGXeSqdtehGddMZ+Sub80qYy0dn8Cob1t75e7mAIA//oEMzNr9AQg1hFh
Gcutwls4z8o4xGTtD2Hhpt3cnsGj9bGMzM9pbZjj2Zkv3Hvz1rBvA1UwDELYoRPZ3jTn66N+r1EH
e7n/qS2Meo8l5TpFU6un9r3M5tiey338ChaLJEyZjjMBE5APUaiomHCxsUwuuOTLwX/Jtjf6YAor
DRY3Skp7zZryL+i106OfP6FfiSHzahnwBTh5LBH2uxwxkaWi2czos+xnebqUK1bDmtNmMN62MJHp
+rshYcLT6uyGCy8EaDb+NOcBf0u9ean8vKzvpnR202iPtlaq+4Q67eRXF0XV+wec40wg4Mobs3lL
Ei3bUgGZ+mGGSSd71wjCaiSxxVC6widwur7asaLzl//xIo6vawsm+IaAN0uLg0FS6Cp8tr9WgMlc
3tDG7xubbYET/5tKk/ZEDbGWTKkVgZuPLm7tKfeEiKJl18KMeIXXStnjNikYtN+Zb2yeR73jQ2wC
O9whlLCrRmGF9ekOleYkWqv+MBxFEU+qcduRwfnsVSg+rNre1qtXYZlppdBr09YzUpqPxnBRu3f+
uC1qXZhEC9IF4VuAcy0ADzUY4T4MoIfZ/FrG+RcTwWzfSlL+JUciWnBmdaCeI9QDckTByWeQbyuG
wqMu6w5Viw5do+qwwGuGr7SSNuYQq2rzJcw++HhUEKaITgJSAotwbDarb6F++2RMhfXEJx5E57Si
AwmADY2uBZbrZb72j+T+/nRCtYpXIec2W5wYop8bt0f6IXTaZnAoMTsReKtPojzRyBJiAXm2+rHN
TcLD2TUH4h5xgh0/7bmIeNJ9CWSwEFm3C9O5JU2jv/9gU6EeURMhIEIvYIig+0Iz2FgCL6LetLD6
Wh29q82MAQ9tkq+Cw73Of2F9hJd7anaka77Zl54ET/0P4rva9C/CwR1WHcRze7LQTfoFBu4lwa1t
fo28NYqe9qUkjGnaUvYU1w5EZ/8+gqpE2eokdoPRU5KDgxfm2TG8mKKxnuXZ5igu7PWA3aizc8r6
ocQw3PIH/xEtSSGEMcHr5wose/PTejy7XS8DWaBHh0I2RSF0AjzV7DJlg6MNkgF+GSaH5w+rL/RP
G6HhuSvnt/BVGJwW9A+NT7YBIoBUk1+PsU7X/KgdtWzdbyg1PqV0bNV8m79UsT2aEXuxe5Afuuzb
vfR9zEac5AZ8h9lt3D7BbAlMqCho7dNg7evvLME53GGo2NHZcE4oDUZBuRryUDp8knhx7S3oIt6b
S0sUqzlinV6SGKLBDxOlbatc9JCPBsUnDhtbwOVCxkgP6U9vPoTVbnOstK8jGG0tWXXHa15DLLL5
aQbEFt4Gq9KRw6746iWd8dQa4wao02gdS+r6wq5uNwol01SaoU/B07j08MOKkdVQ7GLTb7xgH1nc
AeaID3k5qXvlEB1sKAIyNMmBdV4sEN9q84tiN79GZFK7WvkVlNQndubWFNo0Ab4x+2YF2D0Ga9ve
R3EF2U+AFZhGphFLeB8pm4dKTz+mPDycfXj7Gqmu4ZVx/eIKiG2P00Mr2mPQa7XMLNAgOnKCih6L
J1UDlILNQiGZBataHgQQ+Fgdplja2xDOZvnBMf44X4AGUd3VtKzhQZHV9sVwcNCXqAxTt2p7pzkJ
9t30ArTKZR0plnfa1dpA0AUdxDVO3Cq9u3q7dCCm8K9yuqylBfNNrW3IfligQKalDxeoB+xWtKm3
2RULtLZepi3Yi1cWX8on9ooepWX/eSucfeUv1TR5XyvZKvI393xvPBKbvX/ipUY/1mGw2V+ozdtH
Un9iuGFxSZCFkKNbHKA9RXaDwr5kSa4kwtvxfd5o0q7HcnYAEggds1sJ2LJV6agP6wr7ouQ9vnAR
ywdi3YmJfJgJYm4JHxbuCAhstb83VF4HWdFmZpdczcgOQgS9t1wkpZCW2ue/ixoU1No1fYHJnlIL
PRIQQzGUkhLTCtJ+1JQr91bZgjZYvYK2z5i2yIXvXFsXB6zSqVoC7aMF6k33c9JfLoGzcoDuec3/
PO4HZ5sZKbkBcEYQufFfmE799CnvUfG5yTdFopSS5U93Kg9zSznzyBXebjwMs106OsKmF0Ih2Hm6
STD1Y9iFL19WaixQR1Zocq7lhIbiCleu8pmVvlhntc8aeR0CYKBva5F9I0SN/B5t5hkGOKOOAVtI
xPoXH4TcgsZPQ58iGq4hr6kqLrRgDF1m18EzKH92IG6ia+E4x7RIxTcyiSUmmvZCw32blxH+ap+j
ypbCbhCbwbWi7JvT9ZQVUuaTiixiIliAosJJTPhWJGWPkH4waIWKkJZRzSnOODvUr605/SYVY3IB
SnlXzlByqmwG9ibMFSLBTqN8CByQdCUWzyYxi+yY7JO1eA5PslZTl//4Bph3BhgtHN3qq+n5NDOc
jrUyZiXfI/gtVYg1+poX7YD1WFUNiYs9gBGKo7g1nam7Og7N980xyx6aUslVf6R9sA0LHI1m5CMm
VwgYSycu5vc533lKG0shs6xAi+npmjH42LS4XySCv8qgEZKRPPqZ4YZXmUDfoUckBSlynmBzgRCT
XCtP+MKsHoQ9H+MYdsl+rpa+VR1Kp3gtxthJqcZ1865GsqD2HgSj6tjTajHXCrN+dcHFyp0Ampdo
tHKrlDyQH0R2U4uKi0MnzJazSjVVcYxzuybMNFngtjPJ2qnKotHX2CnWJG5lXHdodPoqKFaJJVfO
GNZ4W2Q+KZDezF94w0jRYb4KpF6zm2MEgOtB8NJZAgWDePQF1IZwtpTwhydttBUWysMz1gGQ4jlF
s6GHVkqJDcLxHcWmJHnFLhrc8rYfZFUTgp8mYaNYbcRTn5LyF1QfQjC092D//pV5qvxl2SvQOlUW
mtlg31D1inY8323Jr0h3cXSKpCVcoLAzfBfJ8XV1kQeb3xFzaEvynWMzBcDbGjN0AYsSphgHnHTq
IvRnXw9qnXGphYyGHZCq30TAtkllCbOqQB+nYGjPzKfyaB11ERdj6xMkdqv6juHNgsxrHq0boY0s
lU/mmhrW7q2/thbyiVwW2iDhso2+YJTMNPk9rWtP2PLjQmRKmOk9B5NGR3BGGiTZgYyQ/nC1cBgW
hHfb4vi3+LkSwLh6WInD2cuhyYlw1LKJZ+ayrURCAvX3vOiU8e9fAmhebz95m970vcoIXj9l9wEW
FKDk9gLqtMYbDKa94Il6aG1ps4hEbiYAry9r8vYOqFIM4zTGNpa2buTE2MPOm7ZfdGTeZ851rdwo
/3uZ1qsusmDZja59IkVJnaHmad+MxT1/xYTNZ7XEJO3iJ5iesP3QImiYsdMcK11wenZHNLMY68v6
XH3WJ2fe3DE+vZjC7B4ro10rCG3o04dSjJDzdb2eGFqmMWuxFfNV621kF+Q3IKJ2sPVGd0a1Szq9
oHVI6XfgF6LRfkTuZjo8Gex/oPkLFS/vwtLEOiedhHZoH/5o36LvM0xyxFNwI7qXDJT0R5yAbUn5
sUcJDwFPsMAGOvAShZs4kAEWxMdsYHQWnkJLaotWa87JA1Ru8hRzoT17SDt3LxTnvaoI281vWoIk
k2oNbo9LbPuj6k6PuUiiB8ptuBaoHz4yiZL0CoQ5/LfTFVEcN4viAiSY9m1TR9xXInc6wjwVTeMD
JSTGrPvIxGCtT3wrqQx0dd8P7RQllA1WdKOgII/am0t5uL3E5wnApdvL/0YdmN7O6Mq6PD1Y0alk
CbRnAz5nx47LMZ6RcmmyOJsuGAVpeov2UkwJDSIGBLnR/LahQkbr/VaoN5uplDSCoZoQQsIKzpQP
kmy1eniH45zHKTYFXGAsJBcE0LJmxOgeUbGZtGgrJxv3tTjqm1Cwa9kSqcd5FXS1fWwDy0N4EYye
dnQYze1qaIoHZmLjuqZ+LNPDUzQOi3mc1EuKUxtst7YonTKJcMNt3eabzEw0cuig40brVaT78GPO
0AE7xWIADciQwKd03s6qsMqabRux55hkkbD6+/+A1Sy7c5MeoU+kayz/tOsVlVV2ouEwZNi3v0OM
OQ/qAok4lwyc8D5fmK/yz7+Nru6hX7Y4pAiuLTtmohBLB3U9+WKthjqBlzp4U31aS3uevN0ulUJ9
NHLtMTEJG+Alx/lpbSXsZ9qhddI/E7LbUpyGJmZr8G/tpHWVss+MzRvqW8haPquz5jbJej9O80/H
FUpnXuKepATc+i5sEu53ku9L9m0YTufVnUG19j2WqO0BcEfdbSpZGT7MpG5xBRoNer3P1Jh3mbi2
h+X87ANEkfTR8oisHspB5BlMfv3ZyjNQgPzUF7/4fAC9hMktjIanrffOaWScQOrwGXQSPW+mnPdl
2lW6nvLr/Ry9y7sHtRy2LN+qjy7Inm52JgTFqEDrw25L+dlOAepeW7D4aiR47Ga8PEZlWEhMe+J2
dLuqIOb1tHsvgfZiLPV3SQVeeHFNP9mY9y9lMBF4xhWzKOrmPZaZL8cZZAHkn7zYi1bbW4f/awRN
MTyvrkX1oI/WR8vKEYvcvJlxb3tm5tJc+9auTqfMjGHdUPSV+l2lVBqdG4dPT29uRW+au5VNClpY
9ihZg2lm9HCYWOWd1r+GfMvwD9b//1q0146JFGUTKeXFXazZ3yeH3teOGHwV9w8RTFf9HO1flkeK
aaUg2XBF1DSbB0qb6gGy8DGHiyXzsQdWwdrnH7lN3BCzUGGtVFYGNu470PImw/Liiffnts5XJMHQ
h5XoGbwTl2cA9LCj9Vze4VTrYIiyN4Wgvc22e5P0wrsGvz10mf4z7dEBG4Vq55B+z4/aXvuSBCfo
EXOkP5yGX/WqYC3keXsDs9pFQcD6DYgz6b+aLLEtY9MSt2ozSS2rSg76LCthjwmc+me2RDfL5Alb
rVxGKa02myQamhEmhHOJpI7RmpI01WHUz0ePv9Cy/y+WYb4N75heX60wyX0d81VSW9132FEaRh++
FHP2MLA0Yu0nWtwUQULViWsEM1sek3RpaHxuZqgOhjXW5MQU06A6SnTaJmM+AUdJZcIZInyrrktx
3CUsWj92Vxu+V453xs0w1IYACnr5hzm8Rniy2VsO0r2aPF+M52F7XOFF9vtlaWh6cMqhQY6W8zvN
TbHpzXQjxcNNg8nulws3kc9ae2XC7r/c7YrwrOGZ9ngHT7q7qsV0B1GH17djJ9Wzf0+oKZ1baw7l
Z5HzrqEW66VqdCAtA4JNbqflO7LolfOv1+3jqaK2QbZGfHog2yMh2MuWnOnWcVMnQVTAPV8smJou
CW2Yv5mVNvMAaNRtodKJPTyg78SLZNlPAOUNyAljcw9ZBbMVeK8JmUmXZebsORQzrdqxtPGDGYY6
VKBUbe6qKqIQS3bicI8Mv1Y8eIreQ6OvBMfMc4KwNqcbV6FWVLpReA5X20rHXygKR96xA8KSBKt5
9lU4imVyWj4TxA546t8YL+DndxtuMRiivJxSf8UbY1OqLNvsdOAPBYNTcOryPbod155jcY8pqUh8
PdvhwnZ6gzmQmx8kpt3Hd99ss+f0ATU9x8RvW7oQ7+rw8f/fLu53eVz+YdUGJsGkD11dID5Iyc5H
gsCfuaMbxc16qzKuAvdr70exPb0vE++rm3//4hnNi8jUWQZlkHnCkXiMznYxQtaxWYnU++VCKspq
Tylh18mKMZZk3HKxsA69cgLqQJGG0pLJ8KLW60MNQL1OEdvVtCyeBihyABF37V3zgOLXN7uadTGl
6tjjBYfva1EkKwqhR1wZNV1PUN/jfv8tI0W++qXPW0JBZ7tQO3+QlVpxQbqnqeEsyALETNXjCxWq
WZBe6CGA/Kl/l8kCL0XtzYh6Np1fZ+h4pO2l6UP0sy7XnDy5hCxy8xLQng+eYTFOxnfF9NYqY1zB
5c7fEreKkIlb2qglLygqwSWOYT5BH21jNhOcVNtuqa3p+BsoU1G6F2FnyHnAH6Pt0t9orx+xpBS4
B4E/xK3EaeDX7/JBgLFOnbaazHQLw5MVoc60N8u7M/fnmWrsxru0muB7Idnr7Fmrs/vGGL6/521H
mSTHkVOiN+rmsoCfeekQzT+uJumW+eNMRETgkQ1S3rm+wUZrpoNZxWYR9dg4+z0r3ycgC/Avi/Cl
8Wo+Hgdx/cRklR4OG0yk/acMI2+h8StmotNls5DanheQI/dZnvEEH+ykebR4zBK3tVjME9LsNILC
JFvGUwvXa+poicbA/oo3VczNJ6vN/kD9dHjGQrzGvdEK9DooEZRAOn41rCHQ6afduiQe7OH0oC3z
pPm18fdo/pFoOs3rYdyF7Xou5X8d1N4oHa3x2vAxR8e5h1o2LjUxx5QGgwRxlgZb1GMJiukD63wO
gUFoRfsFSpiJ/RUI4nA1SXPEb/pqzrm/Y5G08er09uptdlcvMptN4casaMP7kmDJ3BVcaTtcaA87
69WWPnBDSOjG1Hkg5pcJMxwMMn73cR2u66OJbR3TVeYp7idgUtTmEw/vdMDCVm4NS31Th1ebt+yY
qxMVKBjIh8yrV5eVP10kTUrUvW8nUahK121XY/Hi9Iiox9ZP2lhB5br69UQvgAstEr21WK1pgp71
Gl57ViWrC49KCn6SVtBFOqUear6AjZit0m8hWheQ/pzoE5Ux7MkXatBCwvAz3I2xOquQH2ButXkr
vOahIr68IubJWCZwQ64fGixE/AFxXYP5bg6FXs6TMigwa2eebWj9SPXxwWfV9XMbn2OPRtatb5Jj
DTsRX8qOWhhR96zRPAkhXHuTgM15WGTxLfD+0u2qw3yzmZovKVnvH6qJk3LLiQEbhFsqLzZTAU1O
FSmF2AF2pX8SJWj9sCi9yObkldRTli2G8BCyLMjkxv+iH7mjlBIFfnhE/oELWvUVZwXauTyeXe8w
uo7bbEXTSCHSnATzSND4O8v/05d0WMoAU897EYdbfUcZaeAYHY7gOJP5OdHKl+tVlKDpcAXhg75D
69BMCfLPR0fvIOZWlCU1Imm49NkfEivbOQMSOS8WB9dxIx4Mx7fLQ2kXaEfSwyVpTYdRSaZfd+cy
3tV/saTxOrl7jcVSnenJOudlyrAUbMfoXdr2uHEkYXLwvwZavk0oibu+Hjub6O653YjxFvPv2Fe3
0Xk9HtSSAjQh7BtOVOXc4+wKOUgWWieW45GN2efdR2FJD4fW5+kALzh3BUxD98a4mGciUh/vbfgh
TrWBMnbXtDup3jDOyY15r19qS7lHUHDwCMepQePmRCIIhaDvnaWjl8EAx2E8ZjezTM/XbS0aHfuf
URmCDs80UtUQpBLRyH+f0jNX5UyzjZB3e3Mzfer0sHpHM28Q0+tBQSfKYpsNI0yJuFPPR/GjniWx
30VWgGx7HHA/yWH/VtMI1cEO81NvxI+deim1kPs3nY9GevGwfuhrmEU/wA3XfjAkEC/3Tl+JahPk
aamjHPDSIYth4rt8PXQnhiYSUKDyBGPpf2Wz/m6JhpJhHo1sUg1Fy6EOGRgu9cDUPdwBC5w7mcyT
Eqm9LhM0CJEyTna8aJXwoOz3hz1CJz3uC1HlbowOdjQ+sWzpnzZn3LC+vjya+E2HsezVuKBTu8qM
td331zfTAsEmy64kgZefWH3cfXZHVQnlLY9oOuddnq8/wGJqn/9BR4ZpSV9tGgfsJBR88lBVpsn2
d6AOq3KRLd+J1gkvg38XHc040kMjbzDSXJlXMHfEtqh3PaUdlTCBNVCShmcFxo8pMQorlMJHUOj+
mvyIsg1Na1Vewt85miH3FUxlTSUi/CD1Lx3ATUPZYR+WHa7jchHXNFfw2kN75gimEOs8V3PfazB5
TiyXFUG6WpVasBCevzXCi0tfMhhWR02YjB415WOM1gXAxtX9duOWOEG+O5NXNl9dQF21KXiiYIxG
FCOGLKJJx1R6QxD4Po6YhUR+/my2YSBQ5G9JXz7KqdYO6X/F8ooFkPIjFIU1sCyaADvMWhhCAYtm
kSybo/D0R2pdPPOyJoZC/g2dt//pkCbz1CLCYWEXKVHP4jjbJOQxdhiaV9lkvaPjO0ydRhoQcvn0
iJDQ4IaCPXsJCb8v5Ff6TDhw87kbyd6KLxPLqQavurTiWjHBuNLz0s7V2amgbVBNno2Bvz2mNWyX
bPiIgq8SDqZBzC1ITGrE1J7/uHg3YrEVL6eqHqRkjeajc7Fh2kAJ+RA722le36fQJ6DlMeAuBlJ4
y/eNDJzpdg5QWVlASmnaOHKH8Ksizy9ZNfiwgpg+uUwqxIX2+QZn0HkAMF8iz+DN9meIxEQz4a53
iLKEU8pr46zCi85IKhqL2t96nF6aqoUNDJp3XZb1DMERILF12xUO2+iEFzxrE1RJcKfsuPN9OYL4
IT+OETGyUtzSbanxdNrnBYt/e1HR6wIf7OemIb0Iabi8VrAhbGZU8EK8ZdTU2g6ma82r1b4W+CR2
Smfztfjyr5Wl7O42GunPZVY5tU2jeg4OGYqeOl5N2SIQnR2V1Mn159vqcSfr3PYf4OwoFeRhjbrG
ptYvsUfuCbIXEPyXox7guFSmB3U2CWGkhLOySWhx436YS6BorZ76mXdv3INSX8YPklw8CJoJXUce
FTUnImth09Wdn7r/JXvfwvxgqSe41/05zUT0+p0+uX2FhTpMXqQjXpaYFSuclyX4qxuBCiJI8b8n
Ki9kNYcnBdxKZ1UVwiFgJDScfCnFdafTMfwU/LfVS9DHR2k63VlaTkbQZJ2X+nf40TFpK14w2GLM
K4knfMs/83S9fb9vp/IurpPQI9G/MbzcuPz6lR892hN8Z5MCTGSw9cuMjIY6sPiLJ7lXKQADWCAX
yE1ppJ/HGiCpsFY/Fyonf3fYd8j9w9bOjv1JNtWGk3odSLNDc8WKUnRqJINqmZ4JyjARLPzWF1sH
Zjhbpp2Dt6rxGQXDnlh8beThRXFoVxIppwPUdIv8CfxiT2EH6N4KoAak9G5pSp8BY8IA8R50QGyN
ycDjzczjK7ztm3B70ZAGRNTurziPtzNZu32n5YQhV28dmn47AXO8drKtPKBhWfddsdUmLp6s353a
2NZJyC/DI0fq0Nk//Alfm16jb3ZxDqK8VUqAaLR3rXbgckvGZQyGk2cSxfgxbjsCsAt3jdKTUjbd
y6jnct8jiwAG3Mfy4E63KIMaUtD+pso4T582Y73FgkAXjSk2Ougw9BBLgvvZVADWKCqXka6xxRM7
KtT3C8KfAnS4y+LLSYefLrz63nofZTVwlMnU+M6izIzbkV8GgNFz5I6jSG5RUHsM6fhvAh2cBAqj
zt1h5rAPmRRNPhU1bfrEg47/ShhpmXNtMmoJrecrmqSg+FJda435lO9bvpj0OulkRu0FxBkkc7XU
CwzmV5DjMz2lksOMtc75LvGUSzmVCwlkKSTrozHGdEH1M4Yge8gE6jHaM0Znt8APhx40Xs/Y4FIR
LRQruwjKaJ4D7f2EpdfMdOva9bG25quR2H7JuJrW2j80JH9Z+9by6ztTkkN8/8BqvhnrrvW11gtd
ptR0Ux5X/y230Y8Vx7YaS/8I+tWoZ+NXFRoI7osjvlte0NEyG/gINbznukxL01Kv4emHGyZtaxFd
V0/nXY4695vf0Z8o0fj/LEXWbMDGbuvudu8A1+Gb5pPs+z/wdkizacL/CRFRDTJkpjZ5Bdv0a0/c
X6Gp/a7W4Pj7J2gQUzs82+ujrNQpVAzmWPcRzb5pq7UF+1vC+uByCLfjoiXckounQq0odnCzajs2
woTWVZkiuZu0ncP4F7dD+bSuBOVLmGjoNo81qq3XPRoQMeTDKdUau6nkbApPUb57cBlYz2Z/JfPK
bHEi766JqH+kbPX1ArEjvaMlvcM6tRXLherbi1/farYddrDrosArPEM7M4SHTJvH/E7gHNXNMY3a
23OrcN0SeWx1PAvH+ju03XGK4dkYnRbi4Pir/rB64SCwrXq/n/Zx9yGUezriMR2SUr1/WaWkT2/y
jIOMDXdMn45VIaOAS9su7BbN1N6ScKOVF7JeW9klN7dbqxgJ4W15r2kjiaz2h8/yZqbeVBrTqMBr
9qId/uTN30jx3B0TOQX1yQj0adxkmpJH9lfT32IVu/2fmjRRjHUqjTbWPCzbuCiPw6e86yph7Lvd
4CWNXCfXHehNuTsIxnTlekj+sh6K5k4ENfXaepfnTUiu0Av3aqddI/mCqiFzfr6LcdlDL10g1oba
0QUIpIvOst8k/zmBkw+rLNQdg/XPLTW7xZIZtzpiQYjZIUUKJGrXUvtnAEyWvUsmmXqVeQ6kaqgv
UZb2mz1D/SPo8YRVrDOa8L6w0qmPfmesyR2ZZx1izEbwTdHM+jj9rVPc+9exgevUj18GI7ZHg4TM
6iEdbQdjAe5yYWRFlsStGTkTM69o6lLMyAH50APYN3ifc+XkrRZmCMotUq+OUJrsMV23jIvYbPur
CRYGYLXSCHA4XYjKNAzNoHQYhw+HYezncrKo25JcKr3lEOYII9LD2HuF+kKbwyEYzE7ZntXoo6Qb
4qKoW3iWUKZ/8vP88ehoqWM3+/3n3vNjV+yCCaTi38Z4/tDxpObcdb4sx+JsUPpFFEP8fAJF1XSn
W/kTpkk1jYaeAAMH5v0l6Ifk8RWeFDGgP2dhgfZTPYjJJXfKVpoLWnvMvMXgkPosOrsU4HdvkL2i
P1KHJjstGmqcsaEqsAVCdQ1DY6GJ+JJrKzs6j/da7/RBMXL9BpEn6KQbgxvuL4bMQ7OYDmnk4Giq
8gaq1GSwOdji++AL3BfXMy5mo//GSK+/4WDwiCw4AjSD74s22XE2X2PxAO7V34KaSnRTUeeJI8L8
qjPoz0fQIRAGC6wUJVQ3e30Nx0cXqmhKsjxFQbORC7aNcOP91Na8D3pqe6+Wzuxre3WZXwt+8Mv7
uL8XvHN/7hW8AOTBwE1A/WnEbo6Ci/fn7HLUWr8W9rL2wh2IU2QpvssRbIYV5UjV65Aad9W3Tnat
PSzwtqFfLmLJk3nwoJHindkUhzMKbcsitYGYBwkiW3hiVvYTndiiHk5ZzVOS9B6dlw9SxD8fHSwm
rpJXKJzYey+jSLpQ4YPwJEumHO35nRgxfikuyrApJ3Hm1FlLoqKFSoFcxIAr3vwxmfGWYYSxwtr+
IDaaMZmMz2Llzcd6zsN3TySVC1qiaAwdQgilKDDSHOKYVRqGRe21B3ueEc2CB+VBIeC3mEI8253E
dcWj19ZQhzmO1jN+62gG0+v0RNZ0nPXJiYe0xAt+m3yrQgQLLi8R97TyspXFBy73UjsUgPok8lHn
qDObxLUEUDqLybprKJkHNCSYm1Un98ug5ObNMz2i/zKatZdndttJGstDLfJyYUp7z6871On3No6l
a0IZYR4Jx9RK1/QA9CYtdyS/W5xdErTUfmCL5DrAY3BChDy5QBgezgwTyj3OnvRalRvSiWDXqMpe
QLbrVAXRq1vEDf8OIAtfdUeJi7O8TkyWMer2xwZqYPrks+tNa/uk7rTL8yCfFHDRzBl0c4lYizDV
apITNzL6hAkKSnJqIlOvMyYP8sZJzNKYFPZEX3T2pflofGHGngRpXxhx28WWVfOIhHyKvcTSxFN9
cx0UV935uWKv6pH8u0nti7sJXzss9hDfoEvnUiiWuCqZKJasHDChDYs6eowNUgZs16lIxrFQ5xKx
LHqTMskXikMl1+RRUvZTqAo5Do0zPMBwHpvzXZ/FM9m8cycz8GbNPC8GPwCH4n0DqM7hWjxxWIF0
0S1E7XNwnWjeWqKACFNgJW8yKcNWb6qQfLW31llQdLD3ESnNEMm91Y/UaQaH6CfjhV8h/kMOMZQK
R3AJow10D5KrnFMQdKrCudnVulyNi6a08TjOfzqQIJs94EQJo+dejrF0bT8+DBMvYizZWDEh2HIp
W0rmFAiKpaoicoG8Lh08K/SnIeLC8ReXf3j/cX/xmp+kUN7U+6Tmve3QjcTN9bNJZeVhx4H8YKlG
U0XWy4zZc78aKg89YCKjOGQKyKs6eYyLM2BDJPpenDFG0aUl49+UB1rkL6LwDtOTrmbxwoHmMhCZ
kNogqD5lWRhtcfywUriZb3GIwKUDVyxu8NjvzviFAA4vfogimTCHCycCgVJ02HdblWtIF5PQ/mcn
aHWIMc0ZtdXQFSbsEWOu8YQArvrcHclkivSejqfelV7NTzDuA4UkC7Jwv3UYOMFuEVV27T9/hAm4
YugRDFeStAp9OJBdVC4kHjDApEXXHjgtwUD1jBQUYCDDbQQWvHl1OrlvEjLU9Rio7yp3GY2pmG6E
+p0wmdAaOeSOYu7Bno3uzeA+sqE/OVwk8KS70u3fDT9olakXNgXXtdD19OwbToNx88LCcGw8vxOd
VKSwRNATICNTgifqFdMvujMW3RMk+za4t0zYhmbvp8dQOmlx1n0zRPnZ+MBYXJtYW9iIJ0b4DSS0
qdmax6zqRGh8WM8eKUc1B8PLOI8MwoYVzwNHH7cMZbwdOs2UV2ZOVK645Aze58HjlVGRYTsyGdLc
PhgT/9iiwZtpGSFwkpfjCdORvYDb+uNYrcpRYhzmSE28H0ZfJzTMqKLBpG7LGyNe5suFQyTTff8A
rayFJigzPAgGf9Jk8UZQ9agqMl9zX4PqJeLq6joCiCG/wG9uTA40awcvvwVxuGxOu2FVR9+i2Qz8
C7aZOSTubDs/OZW22JbpuMXB9OB9fh0Hmy08I2Dq2rbkXEhv3PyRoyyCJsmEoZ8xnLur/+7Y6MKH
Qw+jgyt2iRGmZ0pv0K+yMRVG899Od+jUuJ++SBcS0NdX3SrYMKTqJ9ytwOvkE+Ew5v2bdqJlYViM
aagLsnmyroQ22Vc0omDrXHl3ElP/KZbZLSB6gBPpqo/FW0iI/tpUH+9kVgE4Rv9Xk3n5wR71oVBD
onvrT+GB6CGzBqxUbsvNHmq3JawRlh535RNrFr7i9ToKgFSFup8zyHqUDejQYnjBcQecuCqacMN2
sfzudM0i4Dq25IRo7G31oed/o9orvLTSt5tBqHTvcWOC13e2apRZ0MwIbBSKR2q4kAuinRpz/r9V
3ay/8/b5rEneMwW1VBZWlV3qIdsSaUjG4nkQ+Oe1TyiQZLkVaEf1ED0pFigJaP7pxlJmLhr4WJaU
XbB1KtsuIOBWUIAEY7S9ve9fxxCoy8BfoQ/101lG8UQH0Z8miXgwzuraYd2ScbogSHyutaSAvZmW
YCiYNiX3/9TEnh3EQi00Tjgh/630PWrm+RXtFKUHbsWfb4AIKUGeuSO2jfF3dGDM5E0YkVJu5tdP
gcRDWkvmWKiA7e8oISCtljvi82hg2p7o62/h2MAf/LFmroXD0iw5F9bTaOqtJSOIPIg6iITjzCyk
PoHgqFEgexKkJn9ZkYSu2hOfoTXcTrx2cc9y/dnlnZ4zK9Dh8u1bIOpGKIGgXcpn7FGkQFOMYLWD
p3hPbc6ibDXdUfvmtx/wG0X4tro+GwycQm09xYF2BcNflf/PcCVGCyObIV6rzzwsNmQH/0XnSWiV
ujazMdYda4t9i8boKxFk9b9imXArBijB4nnjKAX78EAvqKpxuWYzzTJZX86Vsrg7jtCTlhfMUis5
Azlk1AVhHu7Q2BQDoeHYAwOSpC0rhMh8j1gpCZ9ra4qpcFyxp5FCHZY3bofN4k2hJ1nlpKmfqs4L
fKlVA2IvpRPTBBy1xSe4eLgfbnZqYPi5eDiPPFoMmZqQSGpzFKHGfdXnd17U5YAPP1+gfecHu/bW
9noQfkEWrbSK93d8QqulCQ+VPynLyv+yy6twZX7KFGYPYunpG+E8ITHk1tVLrgcM5jGAp0pTLWcp
crj7BtY5mrf8PO4l3rGGTHUY8L8/ksdvWZfvfs8Vaa5jaeqfNz0zwzyLVC/eGR+lECwZJVELe3AJ
d4NGVwr5PlqH+t5riB7eaGDbRhuplsD1Mml5WGPrSRv5humio3mEktyHRnn3sV+Cr3TJG2Q6WyY/
uqUkBdTjFtJ1QldP/RUBklfOxiV1L8TEcJX2ZI7NIo0Q8m1bhPxwjl0aHLesALS1jZsfTGnUOJMj
eQqIJ9vYTUbV7Z/wfm+486LZUOLlaitDzGKTpL21wnPaGu7bnGc6DoKjvUVJ5ehVFyEfm6lEUkc5
ecjeML4c7sDvtYHciLUSDp+ncfqhupAv0jQ4+oY/LkWIwW07vj1HEGvqJRVdaACyevNzn07KdKVU
8bmK412FyB7waGgz1o4ZQlgziM1Iki3Y0yia7e2SYWa/IaOjfbDs24SsBcJG1K/INAQvPIBEMqn2
/oHuR7ra2BQxhVXP7oHACFSRmlpyLcS3pJc1/tL1WKprXY9IK8emnJi27o99PKb8uTM1YE7JAhzt
VwnOuZCn8tnlCyMsCrd69+mcJ33bzTVI67nOGSzuTfRmRJVjWWCaa/UT6dpon0FOtyP7SOKI5RWW
oYdBUHnNQz98jIwDkQLsx1m7mqwPGtLD0o6UgFnyYEptmd+7GVHTUZ4q9JqCbdAO4diET1+vxLvb
Q7cOsLOZ+QAhpm4DDK8Y3zdRMnDEn8TUubP83l97XUU+WjbhGfKx52LQtVnLGm0THsgpb5zFWBup
GB25l3Q7giqMJdFFEiaSWG4da/rynKb5gQlzs5HpYXg13H77obke9hyWQt218dqAvPTKPaSTswfu
cNv/Cg/hgNMSJiO5/w6cpAuVBj4FEkEcqIXEjkO85nxV+swxK66gA3+yzs+DrLwOw6QJCWJxGwp7
ttVQHC0HfGA5UtPh8E1LGyoW7E5OxH4DhAMzqRtJD5LaxoCovmua6XTChk7us5/NwanG5mNodxeL
2icwt68/QWOd0p70HPI966dRq+Ks+ZwlSImQXQtqhe+OrMjB+GFOz9SQ3o2VoSiuGCxa/wPs4Ib1
Gu3O7L3oqR1zEu10+G7PLJeUmqetnT0DfwV/LFlcncjhT1sFD/4/ZjjiZpC6i48PZr9ETyumqZLr
1QmtaMvHkGjYbz18Mn7RyKFQK3nVQCKEUjM+cy9WfIik2khFCjdXKS0nwtO3KsMHpGaPv0oiuxS8
iUSc4YhcTvzoE4x75WuHKf3BOe7ee+FBtfx1jnrYdMKCfMYLilfxNGqxXpb+AyaiNTFSbn0F/LHh
b/V/KJkjQPhaIO7FnlK3otb7KO4egJYoMrMeFDPk52HaEzydoSiCbSAJ4JQZuLC2Q7FEynqW/57p
xsWtLDgJX/172Q77FGmwRwwY2iZVPRVJhc52ttJcwj9VliGvAyEyW9sMDzO2Hih731SK5628GJ/W
KOAwLd1HoTf+MJ1SDnQNcPtluDoXhaSSp50y+ulfMP5M5+Y2NKHu+hmipQHKtrR2SfpUSXsFY1bW
L6gFi1/8qxG0wflxkYqj9XK7QcjiTj8ZIrLWJay4QWPdi1lgpv5zoguEByXfySQlbeMhSXkOykWo
N5wDBB6OKLCE1DoZH4OiBUNicfsimGLTgngjbNf4YwM/sws7c+0vO52G718FjHGb0hawe6/bXE4m
dzptzhUTG+9lXh+BSkzLedP/Akzjl/0j41i2aq4qB15NHiQULlcY2nYJsYW5SUoOrEwvkNoWxbGo
6yVEZ9XHmxtdkS030cu8GbatsPQJCvHG0aJKz72YE76z+oJVLkiIGIpzUN0pda1B+GdThcfsLas9
Jkvtzvd9JssT2fWwdhHVjWQYuScAdfnRIex4zHJpvcC+uD1zVcf4ZdLpFO5FvtzBjlFCp2x0r3cc
wtJSkXiqB6JkClG23TZbE/OTWPl+A1GAhGRSbVFTfjdkIaGOWPn3YHfR+bsJS8nKEjfZQvxew6Ek
hS9b/ky949LIcOwvTnlz6SCdm/gHkQIm/Iq5eoDhoa+eHbe2kLBysQmLlJJ+W1+aFmkPytTnPc3M
DCRmnzig9bJLVSxq/8Xmiwsnr+KFnoyoRIHH2lR78lpCp5PPjGzEDNPfh9GOrH38pZnCUkQMWdZO
prCib9mWiirWUYovuUEfqV5RAMt7rTV7g4+sUAyla7Gl5mz17xDXFqVsFUHLJIj0An1mOxsiDuiB
uht1SHnYNtC/ZzLigjvQFDgGubN63eAe8+h56qA//KA2m3mmwZdWEFXqaiJB9HJrvvG/NGHG0khF
l4nFfWtLN5o70/XOHX7Ty4QTLquS0h/ys3trQvMXTlmFQeIPTVajU9V5FpcNxQRSn94Kuj7WemFv
rbbk5FWapr3B5JxGZfvDMiO8G3ma4mSghtcX4zXiReX+f1ChTB+ruqngxyFCzsKhULtIhrGs9Z2+
B8drXZNDUjeMgEOdLug8EBMZo1Jva6jcBVA1dFH8037PAokCdi0AvzzjWPWPqF0JOhChIA3r+bDi
5T1nFjt2aLEBcjNtWn/5ZNtkJ3RSoTv4VIysBjbnysfuuCIDKS60LZcwm2PP8NBhUNgXjB/NRmXq
V9Ecx0FqBQSahU8ITx4u5R9D5lIMw9yWZsjScE3duWCxM3G1k2OnaP1wq0sU3WPjFVrVglPVf2RQ
bu9zNjssqyRIChANegh9iv6YpdtXQkP1OIrlWk1wRuxNMS/v956MqHoFa5L7wU5kNEUKBTkriK3K
3rZBKYPeyhwwayD5qSYtjUwy1mm4tDVCZoow18dwLyOBmqHUqbtgbcHjKd5cPC2R08UPUzENzBw3
4QgHePLMnC9vHUd1jbF4I52VIUeNSBmUlecZvH9yi8x2+QX611rG3N6lYSc8VjU/pz7h+rBDFYoF
qG8F403BuXANtu+lZoIdJnn2m3wcoi3FGcCaIJ2ND6ivc7PcNNPcGIJNWtrYCnoLBdmOa1R9Tx3A
QngeOPAhUxO+nv8IMbWCDSvMxea5n2xIQoaTt8HkGMNqXnahjXq4oVt7kJW06LjClJGTRjwSCULC
T5hzQVK0Fcq1+lWF/J59hJqcPhcshHr4832/MELYq9aDbBSklvcWwp4KN/amZ5/cQqzyk37SNJMK
ptXbvGmd3hIbk/ngYJPiOdUfBXOeF5wZaS+F2YpsLyqfTlf1xh3uS7oRLiJyMvp3OZPGHev1GJyr
Ox+DEsjZMwKLH93zW48yr8w52aefALTYPCeo81GN42KD5mp3DDdNGxqNBhIYK1BeJ0sPvQQp+I+k
+VgX916z5jHj+gtygwlwGs+MyFRBbB+lFFGiGgDQQOTg2V9Za6eJjAG8F5mDtfPaWQDWZzuWqGlf
xcm8DGhA8uP4KhPN40q1aHm/0nrCcyYSHJnkogC0n2CLjIoB7XKjqtc6NTtdnCJlAkZZrfm7B0ch
EVC8TZu2ad2l/f7ImbmPJvs+YpRHJdM7bDAhfuVJqTVHAHZ890kvPvdcdgNR5a4JHKu5dUsRdNqF
LPKPADd7fKbQ1O7f4P5BWv+M1zjul18isgpu5oFaHQGGwKKD4SCbl4Ox5FJFH0riPlXO5cE/KFhP
91xRUkj+jFOBDb//1+lkGUijKLWrkdEVMtS8j6BidM5eocS+zq4CUXOOZgctGfoE5JgIKO6iJ8gf
7okyCABtpUYKc5hOxKNVASA2cUR3QYSvydMeuyRjPqbPJDaTeqolXDD1OztHbvLaZuk/1HZYpXUo
z8rlII/H7+Qe9aIIzN+qYcwDVYOUxPTnzOlXdmUdNA8cwR91AQL1cqd8btcuDYJSij9KOR6gJ+Wv
iq/4/FESFrhC83ynNQz6EH3EKkdaWIYdN3Su7nU6VRPM2anpxVCB0eG65uCZaMFKbQR+SIKulHhz
KTfgaW/A3aaXFvZ0A2dyWEJ9Dy7MGWRqiHlWG8rFUeccvY/OSCzIbbiadavQ0LlyV53/3PWofwXr
A7nGRd0VIMUhP7oZdzxamK3KzvOZRlGeYzc732SQfaPrIFoMcVC1l1wuqfdQYmprZ2YjJGLOQiFp
PSlY1/abxFdM2snNXC2GXlYrH0gJGSGY70hbNVtImFFPSC8JS8LggYpX4Ynj28BHzKHFzbgGRl3P
/6BQ0BNuZgFQliYDujPABHJM4n1UQkAPJbWsK05N+X0tIqyku9Ex/x767XoYa7Fiti4MkYdD3EL1
br255rgiUghbK4ueRvcJNjaM/7Hdr0f8VY6nvprMg7TyK0MFuXLieUnlS6S+hvPvq8c9sjuxx8C/
+61ZCmEm+Up50PhDXk49FlHzK0SvK2ttmKIj4R1Uvc6PsWBjbo97Ayld1W1WyG56lukwvrM/kPkJ
4pMTDJWGx9EunhTuWxffUNZpnmaAwm+J7Poiig8pl7tgAp6aCiMjHTcUopVea7HupZYOytEW9fKF
XKokyR6JIgddK05zIrTb7bCHaUF+i4UOolgc+jZytGYSUqiDpyF+fUVRBsYftFUnyb93G8sG4A6T
KutU3Cn+ZFDVjl5czd0Yi0B2oK3v1VY09Q/+0RCCZaUOOL2vzz246bRVV3vkYYo1RZamQ2jieJ1L
ylXm8HqwT8XXFDsYlEZa7Aclsy0bh2zK11iXrLms5WmEzxX0CF2rpYhhkqpt/mRWoC4AG/d83oIv
tRco5G0pexaJ9PDvny+0mSSYk9ooSENhRAuiOXGGTfTFNdZUmz1ZwWmPyLzQffJCdTM3PGGEbT3h
9cUjk3ieclYsYbMoNVKRh6raWP6SVH5zC2TvHCBSUVzmZek0b1mXA/RoMRAVencYD6Z6C1t0jKXj
UeUuKEOYwIlsKHMcmeh9pa4YxhP1y9fqS5KXoAAMPQdR91zxuPgqlIUdxzR73r4/TYmk4QKZruwC
1KkLLo7woZPrb4sxhWMycMVj2Ym8OXXc1XZwIICu0wiS+zDIGtvnCxMQTZZAgY+Z0hzHb7J/K+oU
dWsA3HQGPno80bs74d8ogPRNQEmbRNQBBuizKJa3I0okUSwm0DFf+gNq/nE+HgfQRBgP7qMVZn4h
SCJ8J/GC55hPF6NLlA2HeuZiyFGcBADIrwWF7Nnc9ncIukBp8yeJwbFj5/iA+VVp7bBBzPWsSksN
YwTVK71A3C1HyXk1cnhAKdoF902nu+/9JgckjGt8EI0J503j/iBFKexiSWBKJFz4R3txvuuj6Jba
65TC6wooidiMaLTO4k9vY+nTo7xcjVhAO1tnMwoIpmt2K2t6GtcDTWE+UR+CfSNEj2bIyQ2BcQo5
8P1Cv0/gsIUgD6OlVy2GdojMbYukBCmhEmoQLcfvvhS0bys3RIRne6Vf7TJodZ8eAmHgUEKoYF2k
XwZbRWc8mbCJX/LTKDd7rPDb9wK2wKC//ejJmUlloJIaRvL4bKUUoNTILhiB8+Vmq6UjH2uI34/p
+yBFwio7+p4rKIN4fPKoKYDYuxosEzO0+krKfixu9xOSj87abJjWBpHFDNbciFc7DSk7ETtHJw7m
r72AXe1eOTMq4lgDsrN3oU6A3Fq4kCov2JXbzlwF/11ekeSAEiZiqlPKBJInmAAjV67N5wxz1uk5
Nm3k9GukmprN3WwGwc9gYAtM5k+ETs0qp7Bf1NS1yDN1crfaZ5yXnZ4TdsbldmUWlixI5rO/+KQI
Jk8AUH3YhWOAj5XwnGd0a7tCelMyhR1UIN7L/lj65Uk3EO6sg6+LZxWnGXNo5ahFLbX4xoVG/vAF
l40XHQflOF5KekPXY1X/8MAQH4+0TSXoooUwac5horTPx2kZEJwtXJ9XRNjCp3v7VrjEEySwoFXg
TsDTUuVblmzIBxgQOJ482B86hz5eDc8woA0ckZk+oh76f162JjPXkFSU+RkBTUreBZcLMJ5rt8/c
KF5udKLcjfXJ/0Wf58cBNLtCAeKcDYXV0YcZfey9D4VGjM8fqxKjSzpKKtqFVaiKQsHUCkrBxGJJ
b1pJuJAe5TGw/MFS4SMEgM3g52KbyehrfuYOegDwjHAzlIoI5UFfzln/JxAc5QSnWUntyjAaFKZ5
PapNQshELVpK9l0H/4OR43SFXqdJy3V6gQ79MFL/9yKgyUiVb2Vo6DZVAgHq5qFrS2NMUa/qkCXw
8ZE7npEh0OhLLY7LFogWPmnpAdLPkAVXRaCD7TTolXucanaoPFZrxetBGSTGyeF8/xwA/9+N9ZRT
0PgNjCJ1yFn2EDBpApPY44HWtLZHJgP43TkRPVSuTrSoi0QB1pGgAIJmvic8JyEQq8HIsb5lFimC
8HU15quQC1svcOzBlTzjBNmnfsRd4JA6K3KpYMhshXOJHn/8qIKKRfR0FtvlNXpZ4Tj0xcaKoRWb
dJtXUUQR9stxIi30JTODjy9cawx8bVtI+bqAbGR2IVzMTheOsoh15NGxHAfSxrfrJZgik4U0CJuJ
64/t3ZMNPZA9x9xKFQjtWe9bTYF0MSGFcnvX5EVBNczQMWCC3AjwhOGFJnrisLW5boYP8RQ9LX/+
xarOy6ed7PkOqdZxiwuBVQ52blOrDkbGU2vhdQqAcghKJYDi7yCIfwp+XDG24I9o2nJutM43ldyz
/wSdh3qDT2fUR2dLlyrvu1PB94kUTp9lCWLvEt3UwSzWZ3Y0Jcg9WW6MGJUrpaVWURTwiep1OaLq
s+ideVRhMqWrbWpCvqXcq5dGLVB2Dkm35f/d7ADu+oWOxcbbeV7ldF/CJdT512Y4K6GfR9QMPKB6
84x5FlGYEnTWZSE4xzCQuyjwVO9N9q0/yNSF4//Q2EVq5sTF50nNnuHWjmlGRc17vQxH57vu/ShO
JHWBKPINmUX2rIQ/ILUKMGpHrmBKMZgMyKPxjjlCGzY9XPxTKkSFzzFTkFXRbqCMFmEFlRbjNw/j
bIfLuokM1/pfyGYhvn+n9FNUWnmkkvpoKV2JyTr4FnsmBb2ItXMXzT2cEDDnmxGvlfXVoq63xcnR
Ly9hhWZMqEveO3fIiU+lDyTTRwsDOVlCJo6IfyTPvXGG31UmmJ+6rBlihsp/J7Z/vaRT8eHgRP4/
BgXM/7r8ghtSllDzqT9uKNalznFuTznSrGYFevLJ3ESFm2pvpeaQ//kt7FcITf/rfUZJ8eFGSUNv
0SHhuoBheY8Oz+xgfoDIkm9XV5nilQFFaZAW16Mb87M0RyCiDAsaVC8oHGOZS8JDsci12LkCwS5w
okUlQbSPJKKgdCoyG7cDjT0XxDusTZnaeA7rK0VSM5MreyFTz+M0pIsEj0DY8u9ecDdrXQ/U//0A
BE749ck2z6hGdYkuUriia1z0grWYCs+h5fcrtyiadsvi+M/DRBvXgpCxDMZEzaQ8Aa8cCdUeDwAl
EZvxwExRACBo48s2tOYo3GK4GGTo6Tu0aD33ONqsIrqRLsnhkExXE7oN/8aqXYEFztfSnrZlCOvV
aSqphAEi1+E89Hs9t1uaq/H3EGPsiYb3IEdkvE5IO35nwg0zeZ02w8v28MkVBUTIq5ltWQ1iRsD8
XWbyuvcWjC9xX0NOv4O1s2KK8oJ38gOLkWeGuTYXEGOrQg8YY1IKOium5aw7kXb47YL4G8NQePX0
8sv4tUg41ez1G4neY5Qfbcdr3b255P7vxyz1nR2JyMlIEyy6NASW0v3cnZal3SdDOuqyfcL/4jAq
pqwbsSUddyCnqIAiG4wIwyr6So/LFXeaIvYa6cqRhqf3PgCBscqc8BrtxvKH1w3uSGd79fJlpAtD
rvVwkyOCPJ//Ca3Lrn7JGp6HBgu1v0S46gNpCbz0iUBNICC2uY98NRx0/j7JVxdsZFKUKKtbw2rx
UlFcuiQCFahecokpc3wH/GriYAZFHMhNdtfKEXDGKYxtqrKBK4tuB/OWnie/+Hwj6JzqoNoqQmhH
dXWcmVT+f273ryPnh8To+E0BkPl4jHzFDkGKSVmNpWxC4GI0vycxrlJr0mjw5qcxWGKXL6HO59JV
jxy0bpmEV+SFlqHVH97Pv1gwpGYOT0N8bK20RkVBdvDM0t4dcIKIQzLyPCxo1cgU31XPPTgmIh/B
amP4c1gZ+b7I9cygEqZafqDnjnyABFs1WdwmPMN1lHaBS6HoH6t8JkSUahKGXclVXc50UKAYqySU
qVEXLMCKze+j4vrxZg25rf+P5mb/nmUaQRQLaZisoybYSiqPGbTzBkKGWLzcll2t/uFB/7zKv0r3
dDLWKET0T4/X5Y5tDVjaMDPtAdZDz5etNO3q+3rR3C9o7+dhhk77FrqQQ3AEVgYOvRYCDqYYTBMp
KIxKV+y1uf92qWTC9VA60HIi9d2Il1WAaxjdJPWltslXo/XR5IHzO6qcdBMjH0SGSGpWp0vqZZQB
BCktXKGSiSMZomqoEFn2L02B2gBULMGQonK/lr896DLzybXBSBB986o9zSN1O/YF45h3s01jeUzF
1f3qUzvSOD8+R8j25mwjgYuMOhPmUOuP/c62m0N/11Ndix62UdON5baEXBSCi55ukyNv9YS6KX+D
3ZYilmMyqlwsOYb82/smpDtnD61hQk4SwgRXz7D+mOIZnjKghv/OtqnBUsdxMEExqLtp2NsbDGeD
aECzIHV1CXIZHYFM7zpr8qXzSDYz0IQmriDkXcB+K/Frww8HK916AuVWy/oghutXGii5LEPlgrmp
JgkYarg1gYSLgxR8Poi+9ZvCg08Qx6iCUR55vxYS381DHJlEDM8donvQiNpyBE6LinTESuep2MWL
m+qTHUv8XMv2R+JWItNwKtfs5x33EjfUsDB4l6te2gQn/MqV54529UX7MG19Fv+Hyzt3uc+dATsf
4DPctPz3+9nsLv1zNAXmtIr+5iZBZwz45YJ8fOKlsfsWbXA4DWRO92QjziY/bW1O6iEVWtWior4W
NmgwCg0Vtcz34dW9yoPkF20ky322OVs9cgFPyE3K7E1qODsBcVUa8z9CeYOTfI8QsOVXa9M6Rq0j
CkgWsHS3N9A6pCWAq55nqVv2e6WIWR5vTyoZurMEjXfcZ3EF2zCOLnFvMO8gV7N4mCzhuXIOllBZ
VbPBwMxNxznhGa3V/LRlZ6HClNJZU/32xvI5wr2NyddhpVRnkWXa6gviB1R16YP3rCYpkq12Iexc
ABPvzDG6MVRpbxxAsgcasINMjuuv6lFlghEztwx3HGw8lgFl9EMhVl19OCGjA9w/tUppko5MJ0ko
PicrP6Xs5O4c7rSBB+6OMLviNv5LXZKtYrYPIYGELy2b4awm/5fFVVEiuKF/yDnR7KYMS0EBgD3h
on9K8wCrbnLMR9x/qE0XM6B53BkSUnmVI8HjObpW3Fgpnxzfi+NEt8NlSywf4CpsZLUkGEhdk/FF
oMiqCZp8vgPSU08t1SoAyNLPIf3PkIL/yTOTc1CmqgKshX3C7a8N5y0wpOv4SbqtTFiqrrTzwt7h
lgkgeGDmQOQCxoNN9uAH9xUwavrTkoolAYM1f9OUV/lOn8+xAZ/L8MhXJ9VhVwrJM2n5zHgVf7j1
XY+zJ424aMm/CkW9pSZ9u7KvT3wcnmks6fGfI15rI1v/YH4CuL3Px28UGmx1tluVTZFor4ze6x95
qh7SjinxMtwSR0KI1fFOi3qbtfvE/ZDxgQ99IoYab233FLrCkvYUmsOmkEWxuV+XkcUoX0MKfLVJ
mOS+F2X5AtWr67Cr8M7XDFhCXF4frRQXu8W4JnqBTwWl8SG2Nf727qvI1TkwP/iCR3xUU9kS0laH
e8hfVe3EVfeZ6BrK1Kt6dTZZRoUn5JgBxvAKu24dXQuXTQoB+xntKTnaSxr+lbe1ct4v4JhOORYa
u2uocs9+pIUWwHKIbEu7JHY68zPCLLcsX2/Ci4Mtv/w3pG870LqaFlQGX6+SjlwMefaoHFFH9uO1
8YjcCHwDSJ9fTnAomKzPmDRDSGjghiN0/gmgj7IO2Rg2IkRtBUfFvyn7m3iSGfjff9vH4zWc6yIL
sRq41BQ+EAGl9wx/i4Kbcr2cHJn5z0zZ9tmuDVGw2/JRUhuOuFPI5A/Gg4HI0n0PpGjCttSS/ltr
0cVCX7jqOD6/wU0tlGEzGzJ0iXvSkXStoL+M7slL4Qmt8fFkQuWF+uJuq8T0KZ8OA310LVq9AQcQ
Qeyr5AvHbqUq9vWp2mDbzWvh3Ff7U68nb5y3opxlLrV8jYIkcsWJZj3F/OV13Ft0QsD8hkL9S0Ly
iDZaCO2ObnfSd8WbdPP4Io2LzREuli8Bx0szI1mnpSv/RotSUieqoqzx1rcBDmTf2g9OQn+QrXtB
gMEQoQnhGAb8QV67CocjvjU4MDr2//CcMde+4QRFLHfsWNLpBXHoKJjL0ixMJma4khLR/vNfQaNe
IwYccjuuXJ1QdjVNseG8ozB/jwlGa5zXqAZCBNVSYr4pNdk9sJM81lGzf0r8AwFOknXDvJu6nNxp
Rdd+2amFz9MPno5K7YAEOsjy4HCrQJyvZ3Mr/qsVyR3Uj37F3T1LvakOeqeiqM1sdlYAoFFwg4Rg
mOMgjSwi4zALpL6FsQeL/Dfx+hxBhvn7AgQCO/u4lywKPfqx7SoZT6xGiCZ665vzoWntSoOoS7XD
S44elBEeOO21l5MjcQVfXjZWHHuzx8jXTeX5MFTVQvsG9XclcPeROQJgupoI/vfwgu6cwpDsrtzw
aCQ03+i4nr53WtZmqib/8Xq40CoRVwRAIhMNT/d6q5MNwiPb9Mv12ab4hvFnml0FFYH83Y+kio6b
iDQZfL7jzvEBKfJtDzK3vGpa5ghGm/JSmtqqH+rOzFiGpX8o7OPCb7NrKzTKdpNblhwQw7tMNRyE
qu41Ck8rY/Re0efHwGp6XzUdlREhm4v4ASu9mbZu9zZ8o6PQNPL6WxOBN6eJiWU4OH0H8IJX6lvW
YoQ0GnSFYrCP7VSSDHag5NvgEP5YEqLUjNAl5ZWXQs3uW7eBrrLKStx7jWwsbZ/ophcRkOlWVoN0
ckhdqVrAk97khC6hWKZxNrAIa1dc9GdtE7LS87pR6ufSyt9Ntcv7xyhoA3j1hao14j2oZN+nWFTp
j+iXFEwbAQEPRFHkeFtrQhgM1HQDeqKuv2a2KiuIH/y3wwvbXGSQFzVzlGzrSJup9Cn7sT4WFY/0
wbFRgPcv5y0OD2+CizcJywGt4OuxkKBj3FRbC9+dtNlB+jVOElubzNm8kP7XFRAA8eiWTT8w4keZ
C072WDlvseH7fdr8UkzfnrCBfQkzjwXJ7Vgrb01GbFucX41HUzQ8pQaeeDkdqd5BDHY5T13pf7xA
HVcNwmwwnpkV+j2ngf170y+akyOSCe84+4BztmviYkYN/P419bfmah9tqX193ElMFtvcctqWVBfP
853WQWEsQIdQG4EYZd5nNuwdxT6GDO+2wjMzQZGcN07F3RHv38C6rTDmeyk6seYcfSjYZsHOG8he
E9LXyjs4Ec9WBfiyEjcnh6Fggdl9cJkPAoO39t9JZPl/A5762vcXtE5UGTEM8m/KnrbOUO2CuiC9
ErQt3IlAFPIsWZH7YzYZPDRPsyqdDpmYrS5BjlexK1wfB3l2lQBKnigtESYluG2+7nGSp6QUA6jn
/Cusog/suXXuvsJWkLRG81ZZB+HlNzuwCX0n1f+7cs/y5srmxQGe3orwEdmEDKMSHU1PXLwq2GZx
kQpjvL16Le54FmfRDYiq8uXD9/AmJlRW/sSBfe1a01UX08V0PL4sSszOmnsEjYBw2wi4xadk1HFh
e8Lz57xhFhB3JGlQCPkqgxW3mP07fqqpgIg4OYqqhBNwxpS4mJj6iH3zsf0lrMDvrY2COerrY0v7
W/63je/SrDhktQ9v7m1UaXXD9OvSA9lB3IdSdwl1Xz+pfPrDnsSbOkamgezebA8IG/n2MzMajKno
xpwSVL1IdhsTW95WNJNHRxPqCnoM6fT146KmIikxSnR+eVijrywB2WCuN9oAuCJ7TeHRLT7NAxdf
n0mgt1fW1tJB9rByzn5pCC46DRd1CbElQ9vw3Enc2dx9Tl9jmfhObZ46s5DHPdueqZ+z5CcSB+zT
DS5edwZ5BL0TOP+U8UA3OnghFDrbgwWkOypWSgMaVxunXmFXbW8A9uiGYnc+DmTrlm0lCWAMti4W
J0EppTT3YiqWfofEYDWIlqD36ECe8PorgWWcG2BSSWs+XGTyYUhjwkhNj1vnb0S2Au8hqsQdOHhY
RUlxZImYKgC0lkEAGpLr6ULADtf8BQ7pf9ME0ZxD47rYqI3JeV+ohBz80Qtpt6yXMitW9y0+WaZK
TcImu05dza29hqSxAHO4hLv8csrjxVvBsfyBMdmjLFnScNsBoA/P3MWNqJPgFUOdrdyNZ2c30gLL
pOzKfiy0gUSV/BzTE1MyvnvhdCyP57oZZFbYwKXap2J75B1L0YwNtIWJfPUafOfkhatwqYfV42n+
PaKXdLGKyWgVuJMw+QdQ4SKwct4kOq5VFziFHbytQZ8ldP9yI1w1wAceVd1K5VmJBFD/HRAx98DV
jB4qIlsjYqZvGnMeanR9T5DQ44z/kZ2NnrLpaRNjlKqGLuQxKNRCdx+3DzLF//VxQQam3hA/zegJ
653e7yxWqidJO1Rni7BghXDWkZT0xmQb3xF9LkbDh4fObs++mBQNJuFsR5oMXCosFxtCzhLyHqLL
nyNTh/dPWYGofm//K2ltxunQrIpKq5+9vlX+iJJbbkzwlHu9iGdMbPJl0AoePxaSPt6OzdO0QDCO
K8ghVkK9+N9Ebw9tIq/FvDOhnE3p0OxkYTJlRnDn9WSZE9HHjHKI5wm+FJbLlCxU1sRuF8hpmrJO
dn3icHHwAZk0lWzdn8neJIWu5yqvmZdi8qzDRT/bHq3+nXiC7BqpmIEeUrPsGc+HQAY+QyYBOaaO
zBZyXn28tWZX3TJNGdKKY7mZoK9TFuvJPvFVMgjI9ZZOhp8FaQpaGNiYLx3qysJhZHfZciSvSEwX
xX3L0slzvUjjwuNHvlq9qctYA92Lx/f3KzraNNVg23cv9xNH1s/Qv8xdTUaUgN3ut82gesctS1kR
nGI4prkUJFNHW38GQipqblTEoFOKMED33YDPvMkeoHIDqrkBn0EWKE7pahwX9oMPFMnSqJgAx8bH
6qNAal0VeHRiYZsmC9rWMZT4OrVPj7qp6ejjsMbcPOTVBNGXre6kvD02xyQApXLjzfh8uUUiIh3B
eECeuWVtyQBOCVVu4fDF7vgKDDu3l911ka/T4Ga9Ojpl4y1FOwd6eb4l5uNZiAxTjQE6sCjDX8yt
25hjpUH8UJoB6FYipF2nvuqWiGi6fA9C1mVYgCMDEBI5rDWxTStS8OW/87vZbc08urUiaBFR9b0I
vgj+iYzdkCMUmt1PlpQRDj0Hl7AeXMcYflpFuqtF68k/Q7xSX5F+K331oO25TtTMKwR2+Fo4lRO4
dE9HyB7HbDA4mqs9+EtqhIWn8Ar0HSNB2AyAzs/tCkUHPooqHX0rnhW/wZc+M8B1To7tYYGcFoDW
yg1Jo0OCv1eMEdXlOjGu6ztxJunbggHhEKCTPihCgHEL2Jgegxj2WKHoZ0nqGLhrql5kIgNfnshm
pGEeP7TddNE1qnaF1HPys9Izj3PjQwp/b/KxPtRnd0BUC3gheL10aoV+V2+bzvGeTTdXZ09hbZoL
CE94J0nqIY0SmxO1ALUtk84exuuRZNfoYRDx/gghpLiyXu6IfQocZ0YEUIyTBNVIM2GDJnO649OX
rnDDuH4eC6zuxon+Z63h50DWnbJ3Wyo70p8hM+EmDDgDKbLFc0D3SaXtxLidi8a1Y00/RAvV6nmw
nYEc8h3Fp5MbiQ48s3yhVul/3iNIo/CIj406cZtCAzTgdcvUwge5uGCJ7sYAeKT3tkEdpiViojoo
pHwZ7rYcVlvm9U8M7gVlPfXJ6fMc7IyLE9kgpGHMFANiXLStgy/c0DtWUtmBXHa1/zv0VzGBJI3D
Wnr3Z2Y2zevX3ekaHMyz+AqmmO85bvy72GhuaJThPJjZu8s8fArWgXEZnkfAPCsfrhbgWltrt378
MPxOpP+gVQ3L2IQ3fhER+WX70qMqmv5bzOOnZ7VEGhuxC/hBYzBiD0x9dgwaZx/1To0E5UG5U3Y7
Qe9VBPpp6uyQ8TrGGEDoRnHS9jtWg5NsBzJb1Ga/v2ryVfQbQ9XwT1X/95YloTiGVS9cYjnCFcPG
bQ4SmCf95i0HFh+fzf/pgZILlbWwK+TosASl/0LBJ8u68MA67Bv/yJ5j9WDP9bUxZs1AeK9pG/mz
EVmMa5J1cpYXT/gKENJLzw8UT7kvAhK4RIeB/TqAiu2/bCsrO0VtBbY/DwXDVuFnVyjwuk9TiRuY
0+oMumhvnWD3iEmHnetNlKIH3HXZ2W/Ze/FfAIaYXhyVWXDZpoM/bgQbAr4xOGQ6D/0zCxARcSs2
cxO9ODJlsX+w9piOZ57GKfV9mOG716Gv184IvfrmRLhHYdQdZ67gV+0YGdslNguhA3B4yVoRFggC
yBL7b+IH3x2mNSTRTrWrt/9Wx9lI8tclHLZRfI4SKYuUovBI/dAu7hWTsEXslpXKaFVqgoKSSp1Z
h0RjNJ4VuAHy8zTNSppQDJYtv+4P7m0IcdYwF66fPw8cykC52zfyIqOeUzb8z/IS524QAuSfwUzV
XlRLrx9xCh1zp4yDHc1LVZYl6LVnhzBg2+aVQgsp5UT0KuXy3QfGT3CtZfY/87mehN2c1WPfIONI
aZnhBgp/v5r7fU68u1uHTQdAhHo/87rlOeESERngD/XoAK1hTVf24G5FVNFsZGSDjPavfHoqFjBD
pFlPBfuKKlsQl6BEwZ7+8R38vY2+yYoY1+LgoEgUU179GX3dJTDrUO7eNmTCFJw99zPYfVZRK/+k
aEREVBiT3ogmhVp3ntol1QQJHu8VVQLtiqALPOU/tpTBw+wUh/vAvxWbmFJRzbKRuD/WA8/pZngN
qIHM5q2fybcPa6gSEV3C3y9jTjiuMto0e6eydFF0atXDHION8F4os9Q0SX/MCWpaHp202EilVuy1
7YSGtMkNN6E3wQA8wwwycDzT3kH1e7G7ias9KmjHzcUpAVHBpffT5n4ffjIuonxwlv8SAAqkNAKY
gMD6KiIMOvWmMYf9Ftjy3ndQ+09G/EWqZEnTT1f+0YD2RIulUkvVZxTli3OOkI0f7P2V1dH1CPS6
WBWJC/Ctn+xsgMP7fxNFFvAQ5fU/fYZuG0pO9vr6dPesHVgxZJs2IAlBXahDQqqh5Oak2v2U6yV3
8h78OB9Xxi1gL8JgyZIxtG21ea1F4HBDNWBPCrk8YUnADXIbnVZE3pRz3OnpPb+kYy13p+DTyGf/
AwGi5Jzg5sYoYPcRh0EfH4RhzP2cQicjTRZZwOWUeBq/p71LlGzUE547cIACMRcSq4d/R7dOEowP
MNMYD9GdfPOMb8yN/vBHwn8afc+cI6amoqI8LiFpW9mhlW8ABjlL7yxDMoNkNLPlLIMnYvOyMw3f
uAoffXS6SKed4+ITJy3a88iorN/GaJbefJuTMEmQWlyYAcBEjw0ROm5XDrTGWOrD6ZCOoCEAwRpR
iln3WzHvK0C55V3lTuZkg5eLZpKBIFPj/3ANxcFOgs5BDRYhBXcyAI6CXJ+xC81YLPJ9ZXnNWJ72
0uIIaJ9o9FmMegcB829qgxCySPKuKuOVTtXpZREtLpRMmj13h9wW44MEl2IohhTfhf0ksmGehtuX
KSZaxBJxM2T55mMyLOKJmj8VMuYa/GgGy9PWL+NpvvNQZ83Dsm48JlQnOiHDwMTcg8BDeFk2SBt6
cjdb8QiMK6iKzhgp+VqzXRQkc1svbxcWJSHczzASZxuf4/7uIKfcMCvYKqZXzsOBBtFbMqDWrshf
Ly3D568XOtM0OdeQfnmJcPw5ozBUyJuFxtZoYoco8n7sUPciIn/8+FA4m/81MCoWCYGInd97rRNZ
PM5wMhCsZKjDZFfALg68pn0HG+5aOf7nswH9MSCbT4ejH77rjS/3x5QawTsf2SVCsUAmtqRAxa47
A/4UohoQITy1S91ue0FFTRH+xO4QBBhsOE/93bU2eUCPm5bMSCfsrbn5VR+RFQ4BtZxXz8BmHQ4S
iLnBSPA7AmlK7ojyOFhR9Jwi93gOb+si8bvNGJvNFrGzyOUrSK8DG6GfPSv42Yl+1xF9TRHkqk4m
+48cEmT9D4gmdIOiXOkgQVtSwXhJFHcLcRza+4GZvF5nY9ySypB5ab2HsIFOhvz3lFEP6/Ov0Q4q
tKEAlO/Wfk81/Y+PTxue4nqJDnB9GtIgy/Dp2fSep6pzkNK6xgR4oUF9uvI6aMVgHyLxCs6ECqN7
Mt6WJRn/GcsU5GVZTO4CAM3Tq7ZzYNtvxowCfuVMI4VWKlKA1rFEzBkmO4R82cE3zqo6ILi9YmPO
XP/t0OWPPnDt4XqAjri00hqm8xCmux7ndzA+bpUhMUFB7tpOYADqEuT6q9xMQ43hm9c3mR70aGka
JE+kygunM4vZer80iKrmhPBV5jcPTEc4vkp6XXbnmAmTvJfyI0oCRU+6fRvdY/2/HPYAkgfSLZv3
VBdsRz28QNg7gSounMpvIwjYJ7/shdb3myEaf0xSo5g/ruvXlGh+EU5E2jq38fXCNA6ZDq/VZLiv
HhXtJsuruMBXnKG5ZNmmauBO1wqrbtEF0WXxLFF2/z3Jt/1Nvd/pBwne/UVo98DQQ7n5MWx9Bvnw
R0kLZ5ZGJkJJpnYkV6dmEEH3knCdu77fNrkYYFPzyCDV+ChIasfp7VTN5ZgYyG9DGdBuri93Mfy0
gEB/jv5ZumFPdA4vLXS6ZlYMSj9IosdPkvgn8jApMCsT4POFLZX4zenFeaEzvcBQsFtIoLTfChYL
ftfoJ6oSaYW18efaQ87tqxskLKhcoqvOxA81rcJyy1k2MvlobhoUQxG5AafH1eV1lwA5gf12Bz9U
GFkeiXo8fsSuMa+r9pVup7dubkMx/+fkZTko2yE1sr/rjEOIHUseSAvFgdbAYwaZjhFosqF9JVoG
k84JnVqD6Vm9apqHVmQeaTkV4QVUt+Z1tSRUdsoumAd3T6fvf+QIEdkPtwxWr8gi85De5VUPkOtn
mDcBtKk7zv31IjlF6h1R3izrffPWtSSg/udWmRBHk7fhOXujE8uVxWQAR6zeuH1CvRQ3oJXzNv41
TLBR7V0520PlXTeHY0MhEVniEjFwm1ZN5aSwi4cA0wleZGuEzL5GNPgTbeLJt5lKzJ3wRZoz77DU
XKV8x3tBLJElbAgsgonUHm4pIkDru1MLiYFa3jrfCqe3038cKCKei/TPsoI53SOXfnzT6ltwMjVl
mxSRVHn0iDlI7EpjA5dyyBm25ciE3w/Vd+3+H0lcehD0Dy0+BLI+r6sh9mChzZvQL6Tx757AzDSw
E145dTr+/r4BEW+g5FrJj/xwW3lI8EGtOD1DgLs6ZVK6EgKG+J34ozP4Y5G6yngD4ND0JkT8kiX3
FskKS1nqhFqThVrPuUXnZWwiVKbR0e9nWnWMxGvYnoJDmuLJ2NAeqJNx2Yn9YIh+UR+Oussa/0FH
gaOUkJOe5WiT0vhyP7ABte+BAU822B1KfmizIJEke836U4RD5OeefHMYTqtkNTYjSA64xY3+Xpp1
LguvBfzd31tP127VPGR8mz4ZlLxHmD1FFfRO+PcYMo7RrXiuaKaeLO42L9MChy1FWpMnAEWEnP5r
B+5Ep9QskWMMvrf5qaGxtdMnlZM2orpuoxI5G5YaO8e5ShwmFkJfo8EI8/xj54IdZqfl6ReYTAGy
Pc5aW8rbXEvTsZW6fkha+p0++4Innl5rzRG+xDTk0BdIZF5YuziOILVd/Gd5wRGw+QuSOnciJfrc
v3Fu1AezGZJiHIkoXzPTlPU3N9XBOlL/0ftf5smeX0gAsOaSry31mMQx0fbnIKJr6NbUKcwOujGH
k70bVuGoGYDlO/xkv4B1tslpnvecdeS3J8ITfbRy2gyssRkCenhrrBqJjnHTsGhFOB3lW6qEWXNT
CGlUMAqFVyNfDhyBMHzP7pxpXKGdslBpt9Jhp+9CcKnAAcZUEuCTzJrpBa7IC5PPNP1LGwSW4w/r
hpf70K+8MVnB4HNNfTPz23S31TVZWv5FQgKmSizWAB7bdFgiU28N4oCPWX2gK+AbT7QfJyqcqE6g
+oakxLzKxXfAFDhZXtt54J4+7U9l9IokrVM+FoPwB7oRCO4e++tsJmTMI/da5qmo8GvjMWMcx8T3
9AoDGYPAb+UrZsTZ1dUOqpHlsnn8O8BXl76y3m0/d+SpAGdr8VSZeVByH+KBL0szJSSNvwwlpFbT
ATwcEhzCxTrL8z665f2quTtRtwneBcPOHs9QhQKsrmFn1bUqJzEDe1J4v2xXmJ30DoY6je2WpG5N
rq8GEzvkdm/uvAWh2fQaeXthtyPK5B6xL9fUonZU3Pjqs6D+4E/5ik6xeorRvVZ7f0Y5V9jaic2l
POzillj0jtC+dJahQaHm2B04cNn7NoPlGopTYxGE/gQjDINus/UcoYlEdt3KI9x+Jo4WwbZRVzNA
I7nQ0CE63AffzYwI1QprnU5xgEdzCkH8Kw4fMt9gT3+Oqy8G4cqbvgTRQugflGz/vA8AaWXMDNZE
OWsi9ERfTYeB8HVAAvPgiT4ZrO/Q57khE9NeCbiv9SCR2MZucmI2y9mqoe7Vc1OTZSetzv/vrF1r
SPbWIf/3B1ppcNJmMXV85QcCjI2vi6hj4EJOu8vamA5JlY2GZdwijo6S832bo1AbjXxCGJrZONhE
dRhCL4xXHh2bJfdaX9LxjjforIFdAisPBcM2XNRhhHUdwXRX6uliopzQ9m90HQoB3YZbXoRBDqe/
yEUu2vAfH8GYWRAFjovQF+cHsEYGyMrZ3ZOHfLazdafQQFeBh3tyrh4HuC6W94b2+fSedK3/LKxi
h31ccrvI94kGs/GHGjIQUOYooLhzjAXv8iaPXRS442Xgaxg5QDQBvdUClhiE1xSxGTJ5ouRpHwlI
bUTuNLEhkKWUWpiDqb7NbDciYDWqt8fOYhYFl3a7zumV+IaVHeBC67IjZJhY1pFBvggZO5I/P2SH
B0uQSkopEWAD6F8XigE0EpDwRMM5zBHSCi70gL7OhrbbbeTyDLY/I0fRxrzLKwBu4qK0cbLmEXEs
dcBenx8AFBJqMoAuepsNJQ5xitoVWpxNOZBQJoEOulhGzX76r5S4W0qnNaxBZOj9qZBO1GcoXOO5
MEJbAO9Uk8TD+PEWqJLLe1Os8uFPB+0T0GthGVF89QlGjgND4k8Uftfj0+oQk4Ko+yk8ndNOrWgB
39atqxp7vU0M8Ss9d4HNFwwhyINl2fBU6CUMzavpxa03E2TnOzqQRvUSHUjV4des2mSyVQVAbZrm
6RvWHZLwKmC3+MpwLg4YPTq9wtrIJOqq2Cc58WhWqV81cuQiHQTwjegjofoCU4FQ8i47EFysajB5
kWDaF4sNHiMtTWh0BzwYDv96AxVoAnE4gr3joZUx6w1GxZM3oezuqCwb7/j5Yy1cLL2N1GdvPCER
ZXVqjt90brLUHJXeciHVSfysxtX2k+6t1g/dlkyhLmv3Npau8/ui/vVFZ3BvPszZ42j8RBYleCZz
TXumz72LirXSpTH1sALNEX3gENWv8yEnI/rLstB6FYHvaorKIwD+6CioDrX3DbvXLMVuS3LlG274
GOFid9vgFVrS2ZQgHT4pAwGhIKt5WvzC1rDC8OKZqz3OkYB+2BMegQdlv+yyENyGixTSOdRN1GNB
evX/ttmwilznQOiYWhI6+fc2+zOPr9qBtf8Hlffx0Nd3sbWJmL/txZ1/zqysNEWZCXfd0MwCSl41
Keh5TQCy+6MW71KRpLWINAdSIrHXSHB+STQUfYISlOXeGfuCVST1Jp7UbHH2Ys4yhi+2Llo7bifp
oA8WbCFf2LiOwHUrC2+u2S+3xRM97d8TZ9FXjEARkVYDdwG4UPCp5juj36vJZslDy81mBJbI17NN
Yc1L6HFESgw9wybYZZZ2yXcpW8NNEzuUVY1jn7AT9jZrt7Lq4Ktj7ztaT31stsAOXzQkxKeT2vON
Bx8h79Q7XgPc4AayWHY51jJoKnJV7EYgCY3nmd/bGU1WOdi9HBVszgGO+azBC9T92xJ/xH+kfFzM
vPhdLHN2SndktnM8WcX+1BKGHfqrXQs0+fhDZE+99f1iXgSsXd45G9b4jf+AakUDqk7uZjX82lb8
zT3I93hCSsASTGCxwFkKXKiwCx3p4KEqQFVZRfR/c6Zjpz7rajoPsHZ7Xkm2jXwQAyQxdjugQnGT
B4Ua++ld/HlKPgMw63e3V/2o/sV91iDTzjxQ3MsmqiC3hcAfqFFjQWSpp0RHAGuQE8XGP+TNRVF+
9VFHpqtZCYvQNGkxE2conEcR/aAdMzIE5Q7LQmBRLkL0MPbELXEy1BWZefko8FFXQiWuwMYO4dR2
I+KELEtESo8jHuCUh78dI/s8BSyG9fUzhpjldEaLQDTLIVz40G7j/kPtuIkmkmt+jI17PO8e5npA
z4dupFB0X3HPayx7SaxTcG//7Cjzfb38JAou2gDypHo//pnBbr56j/L+7xtSiMj1kZhLeCBhEaOU
pBp3P94uP+80Sz6vjQw2qaEFz//VT08/nIouhlGMurMOE0kD17VPISGuUNIBZQLNIILmz92IA2st
XVts6K+iKR2bciGb3F1HfqqcdKxxQ4PXe3/8NTEwFKWwa9G/Wi4cRou5Si6zxCzwjxRs8u0+weSU
5XgkcYbR7eDiDcK8sD16GsWzLqYhtM9sGwmLQoErOTp37X5P//+U0C3P8o4hxjCNoFpzI0aoxx8P
77QUqzS180XNgNbTt9Xo3TdLLkJ5ymbtoS1ocm3f3SratwC+7PGmrTTmx0xWWbXSrBed0pvT7OMK
1LQmKWWUmJrwSRbUrf1+aUSHX8uUYXW12m9WdRi9SM+PGkbi79RhvPrV6OSOMcs0TS8PQm0cLsvN
YVyywQRInk9frINQhSyBK/wDv4UIN0wTG4h45Y+R1CYV0DWd3K8ceLAKJRFNA9g31sal8+/OHPFS
BGQAKl/CZJKMu17Tqpie4PUXRV3d0zeU+6yHQW+KXGGEVmtsPLbQ42J3vRp3MOP7EJnpeOuVvCHS
h5CbuJoQOrGX1A2dnytkV96wysJm61+RkbX6O7EAI8IGU2HQev50uptDmsqiKShjrg0DICVbKnX6
GLznzbIZwCIb3RXErhVv9NHDBeS97fDVJeIuIJc8UBcg9yKrNQW+hB0o5gSB4NBUGNJC1Ef7hH7I
3U4kyOGi3pAa1nnW8zVdg9Lru963gpNGilVOtvBPeePBvX6yybf3XCd+bE9H80CYi1JvgFgYK0IM
oSK+F5rB3bTVVxzVFNwRdejXFzUFOvza2Dyu8sL/oCmaz4wc6D7UhXYTQsWFKIKx5QCCsVjV9Dvx
KHvshGS9SHNtlaF57buKs3+l63yCWZhpU4GDa+etIsVCbLn109q8yalvP2Jo3tnRMOPFqmh22tu9
s/QOQfoC7VSl3MyL4BmXpWkinNYPsxdv2ysEDqDxzBFMc2N3pE5QEVR3QSQ65MKjz0FBufsJlRSQ
tgOfK5z7xaUVI1LzfZKLbuyXr/WsySHRjPg1a4amPxxHeGt99gk5Q22ah9FPUkCx4nkw/I1eZInX
BgbK4HR3pQBoKd9Jx4NduN/2/2Q0SpQq6WKyatXnrlN0aPWjgCI3XIsvdETgtsGgS2ymwAfa29+r
hXNhljj6QbdLRwPTXz9NiEGgPeBx0pLVGU//U+3FhMIYz0u0WfalMtqHzuKny0P1FFqAqdEfLiwS
cBkZjrph7I8pBLFw0jgbVX8V+ytMdv9DfYkBOvzaC4mXLav6mUPPjD8VOIZ1dTZAZesFkdwxbvYh
dnhMAHPYGtMeDdu3cg2VKdcXmi+MEkkPpn6cYXTlLqvuaT8u4FJio7V9hZXdjVbklllMPju1v+qg
+xAdOfWuUWN4d2q/O5kdhamkjH1wmTiCzEQI7M0jLJsiveJdSotsKxwg9z6W33QNK03VS1Lh74p/
h2onnHk4jj7XO8SYeM+3C/HHuq+GoSWSuEo7t5EI5u5naUphx4i8YK5PTCUmhXTroDtwjVSEBF3H
CFj2ssIGVGqWgU2OmnPqq8u3S2RMrQDQrq1fc0e2sGkwibhrS8d8Hl5j/y7AuhyhVALXSPg4amID
VmcPQ6BQXYUvafkycd6o0IO60iBwlYwcNdxtBHwoLtxkrKdatGlNZneJ9Qrf5+sn9k8fARj4b8LH
x8tj6zPV4G8A+RwzhiEBbdXQ7br9hdSVBZpN35fSf6kFwZR5QBzTc+0ZSNy/jJfmWDOI2YloBBdO
WdUOX6EsuaRyZ0ldQm9gyjXhRNoyQpHGSC24RLZPbBb7CJhL2mufT1dpSAtryir7j1tG26KZhPYz
wobvFnSssGZBDonu80SeDGZnIcL9Qci64B4wLU4BCISY881itDUqmI5CbWg5WLuhBf+kg0vNMGxt
NEHBow8tUPInjRKfoZMPZ/4ITZsJhVs3xH4O8a8+VucswyoSjhSKZtgQgVWN5IVAqL6/tAJ00/zA
ZKFq30rTC3eIkaLNU5qXGp8B0SMXADPaQfgTbnJHD7bCG8/Tbjoz1xlIHV1Cl7dWnuKvU67uCHP0
EeBB0H5PUXUXdUvPQZBXp7za19W+jHEZJCnsOAaTaS8Byid3bmq8qpQ+plIh2UzZwaSJIo2pMFDG
MOKZYYkPAEWqillZ4WG2Y9hhRRfXdMmg7J7FISETRKuFxSx0/KH8Rq+jj38FVvxINnzF5jU2zekD
bQ6TzzmQieyiusrsqs5WfZzgdJ3xVvJzVweaLcXJdEwMgyF80a/D9snGqm6Rbl9OnkVwp09+Rf2u
IHAS1la4US4vUZ5TBxf49g+l0dXv0WviAORKiaVpZX/vWo0R4QSz3NzuRBfWZi0TpQq94q7BkPar
/bSUpBW72PK7QTtHlxGwP5HVA/iAZrTBC78r5X4M/ss+qQXqhCaxsWrCfjcIi8ahV/E5S36/FiT4
YGviH9pk1td95qBpWQTYKW68bYj8iZOP+3hXBjK2ZSqhv6hwZW90enFf5wm6jmpAkTDyJgw/zltm
WKP90hWxZqEdHA5PWhkUL+xUn9c2+J7vFdgeItQTLYCEVSTo1RfN1Ku9I5pRXEPyTmy9Xs5HF8Cm
wgSNcOVPrdP6liIspgFUOkygst7pSTLcYf8ReRI4RO17ZADbm6DRYhE+0W+OrT39+VKc5wGtYk4k
zi777b1SaIszv4W6b8dZNxgvLW1xnaywnCKKJOlGujmovY8Rsjga2y1ulXbcsatBvOLbKzVH7MpZ
jgRkOykJiFhzqxISOZeoEjkaD0bG2yj5N7AZbp683hZmpfJMFPUv96IS3lTjtf1bcQ2CXTtU26zX
nVRaGRSMepKVLobkl4dA1/tGGNy9kx78xbtYF2V2vyYl7zCJ5qu0QxHiCnas7mcXaNouEjUMW/VV
VAFZN80XYv9T+a0JTn50xcib8SQqSq6JRizi3V0St7LPktdAN+gaIo99M7QdNwe8BjocB56SbqGg
CBIaIufQaZ5ZEXjF9sjoA4N8FSYhcvpsjcBLnSoTYfXYyy4dA6UYNsyFOmSS2HJ4QECCyes5XUnP
wcG0+93uRhlVYLQn92YWdROmsHlVs0xXyy1vM1dcO+EKKA9zK3Du5xqly6fYLXSIcCYHeeu3Au7W
sYcoXdLC9hLXuyx3ZUYjS/cobF0t8d4aJmBQnhRdT1E1IDaVUznM3cheuBQ3bt9DFcZInuSAl0a+
2PvmbdE3m1lelR/7qh7EL6atK4ylSyCS8/d2qPOX1l8//VA95MbiawTbgQoU/GQjXsVAsdzqhObK
m0svpqo8lVfNc5igmgOlN2Umxh8J+rhgVTXVY+morMylzdr0Y3QcBS982W3cWJgJpIh6r/lW4XBB
wn3G8Xv7MSgWACd/d8a9EAt2yOETdLv4HqBV4jzWpYi02/UVzH4e6VdGOclv4TqHb7mLQxitemQh
1/CCdOsifIaQiqRBGYPftVsScJdAJtAcAoigUwfrkP6E4eFyepCw72Ha+NXs5J+L7tV7imyrBoUG
JGIIusevPnmAK2lAWtvWstptrpYx3XbwIAb8UolE93y3dkDXsN50tw6KA0SBPLgU5mKVrNXyHbVR
nh1tzhd5eOOsVP7nu0eZjCS8jNLHw6OOMcC+oSqbOmZccqoLCNBvaX9e492YX4Da9tY5KC3SwrEQ
7Q0K7PAG6/MbFfvYDWvbsodtcNYS/tOKsJ84xqOduWL0V+fA1bwiqQOQtng4mMhUnrui7F5uII04
mQmHsQB84Dp1wuXb0qIeYCdzUBNYyd4eb2KQ0gfwoYOMFMnK8PgZkkbnnhkLePY7BwvU40k0EeX0
NEbuNhfLfFnb4l8vMswrherHFAmEq7dm892XBsnK2UsE1qgQXdYRIsv8BUQO/Woq2KVVOeGztr+B
XD/d/7aNqPIDp8/cJfsFKpKhsHbXiE1CTEQZKn0A9notmyYkkLilXpk0lz4uS1ioCRvYMhLZGUm0
hEbmQR3buvW2R3MgApNRqY6DAONKmeuMrgczZblsggp5xCp3ph+FXinXN3pvn2PAelOxn+ZxIVqs
rkihrircH/MMOFZqXvN+OV9vE2cHpMisn9E9SuWS7hqUDBKY7LmrBAE4bcGOvcyY/lU376JLKXNP
cY2+wM5kTK5LVzcP17gk2+RwJ9+nQNyiCfpO/rpH11ZYGIIzxcFqYf23riyKGLdb7MlklAHnopY9
DOYNsfR4erQpH+592AvTinQuDd5C0C5KDE+m80RJgzzgxoPi31wEDhrGcOhMs+IZ5qCFi8W+bNzD
j+E58eoeqW6jzEbllRKDayCSkEwa9XWWyoE7ElzxY3iYgrZruCmgCg9NL8dJecnh4l5slfySf39J
DebVTg8rLoQknM78OTp+jzdGZE9iCNRl5vkxrDvD88K0Z3By7EjSlzdW4nT+nFOAdencpv2fJs5J
V9WBgup0PJFXF7fphElB/8XLqaEKyao3I99DI2d9+2M2WxLLoaFwjzvbv6YT42aZSlA57Sypcvjk
lJEXP6iw02adtELsEsOPUeDl7hvcOryqpGnGWS11uzyNP+iozljoJzSPvSW/uLnJsezYS+LGIhPi
lWAqa3fznG0YIcjmjthEy7rK2aDzx/zSImkE8Tj2a1F7CX4KKRzio1LkVYoB8XiduksDB0MdysXI
8OxyF2yqa9SbQMC3bfssv9BZVNpSl+v/6NTor6SqiJQUTVuni7PehUTIFZGr5qyJjQdQmvkOshnD
3yPWzXNlqnYOMFX7vub2PB0rtwwI0fx7479GFdsf+L2ZEpM7qxE3f/O9svEba4rb6pS2NZX0HGmq
cQ5Zz+U2TZlGj1YPicWw8mCgo1kPMjOgbHS1qGN+RQdhSNcVhUKqFrXVrYqasTwbbk0WWLs1K1Fm
Oi+FZ0S/FPuRecbTzz8XHHn0aT7nwEXThWjEJjiWuekzJoART49iF7M+fmyD+8axZI0EBkROlEZt
wVwkdkvJ8LyWjxGx7Lc1C1TC6SMgfKBlsSSA6Ix/AeY9mPG62bs/GQJspZhAkfzoc5JWsefpvOSi
D1oV4uhCJZaYMGu1AA2mt+ZBaEkimzj8TjWBNNE26+rjx/q9rEmzHcWXBDzzDTQnvrpdEspgisUI
mY+GeAzqRFJfSvuUjCZY3kBi8HOMz2gT63+XPFFhq1tSnPXpd3poyBUKs+aIyItxP75XuoCMJ1x3
RM/RQB6eGJbcu+OstE+hdj7dY8B5Qk/zbRKalOSsmDb5TUHUI/47doRYz3dsK3YGUv4p6r+VoezH
1V9IblqmelQSU7InTW4omxYjPsx3e5zySneDGC2D8f3nGj/N0iFsFteVXurt3aD+Jeoc9tjkI9hN
mBmF1Ux7xmqgBaTcgwdAUaPCwxyzCK0Ex9hRLYKatmoWXOfNK1XFTveKWWy80J9Qmsc9pB7bnOq/
k/9AY9qjGntnU1EOYhRCw2mi+j88dOFtHtJtGByEIwslYBb+lFnqc5mFRNVQzMKVhQXIQsEBWOzB
PJQLeDb+ERkjbsBY+5oU3vMp8Ofu5VbrbEIInd2HmmQPraz8ihU+NuFc26LnTtSZD6zMpdiSXF/8
rMeLkUH5kYOBDEeI2xJyVpSRZ6u9UaW9JuQ8OZ70xFo6dgcWVQIaIu3q6keMR4WckqXPD35aEydH
Hkpy2rOHTOY0GvwwChaus03nimkpcETAsIchWVmzj0zmESk2g9iSHF5QC1qbvm6fhuY7gsBmkPkv
E8CCPMxmiw8bMit7kQx2qR6Xf9tpN1uWE2akQtp6B5eUdHNBsYE+ipe4ybEMPVjjboj9H1Pye8j4
fIF4pS98GomZPYfszIvXg3Zb2eH7Oi982QFC6l9QzOxbFtEgV89fHNGVfDDau9Z9x6JuSmlAq/Ta
HN6Cpyl8RqD3gsyrXHsp7VkJQNHauf7JvQsFISr9F0pOsV14CBWmsdV1pEJAthvfZwDvWA4zuPha
xa9t67HAAZjq5HSmdEP7te6znPCNlPagec+Em7jRFT6OA0XbR+Zt571b7AMbTrjuRiDbi3sncPPx
UwE+Ileqj8OXOa44q1QnnK3axcmjiqzKTF8Ed6TP33PJxfcicrql2VMb7H9+OSj4+0b4bMsoumYE
TayZP72GgDwofOzfOIR0Jym5kOrXAEYcCO/R60ILqd14wYqk4k4qaWpVFrmmNFt13ayh9P6WhjXO
urZgQK1zd57Lm8bOw69sMF6ATUkOXQkVstXBWzmnTJ08V77MFoS7g3C6PI34O8nJyUwW00gQsyEC
IJgeSnWn1hdQIxfowL+f5nA8QdZ8zLfZTguZGpccUWIvPlq1+YTKyftqkxN32CwxfwwKKWWp69UB
b/aWcnuEZ6B4kqc+yaP0YTad8hk+acZd52L2FPEnioHASKqgnwCMSLILWHEpwd7NfnOy9D86Qb/Q
tfEq1r6fa/HNM2A3RJ9Qa2eeIkAMnCeEfvZzXMC+YAakTVoidR3eWbUKlAUW3mFKUtLYbE7UjDsk
akdClpp7kdPow5kOIOLHZ8k2affFdZvF0P6rNxXDvNAhLbvnpm+T5XKOJV0oy6g88U5RfUVVR5jQ
fOn1CKiqMx9vLM6mtltpj5Z3ydVJdjzdLKd++KCImUK9v1qEn9OHMLotgyhsWAnc3xaKHUgNuepT
mFH9X1600RnVM6vxncnQpI0df+m8aF6onfon2Y0H/1dx/wPxOeK7ovXg4YOsi/9Omcg2ZMrrD7u4
iMOLUlwsBCkVqMMIvMzE+EluOgV2E1zF125cX1Jht+lqlTY2lVBGit/bT3P8S2NcfulBas2o5VDV
fPH9KsgrKI5ZtpN7zP63+4tQSz6h5GECXUl5gWdQWotwdoMxwCOTRuEST0c81LfeTTYv/zCoL+Dt
ujA/llyMqpFM/11oga7SLmJ7nKwRKnFHLYmkHjA3NA1VSn+CaW/kjjBXFh34muDzK/3jKhxbCR8t
C8fAOukHMB22yGByBLwbcRLyv9MLQCJ1yb0fvmoy5OR+YEcdIZ6DXzN0NVqTFM5fokTx9MNGatqz
+UB/jd9XiBWTSl8d7AINzAuI9o8QX+0IMOmvYUuxmVTXnjqkJVs1XDRX5Q/0utwEQdbqaMyhxw8Y
ifCVSZoN/2Qx6V+4OsoXbZt8xjpXyUvUyuhbUj6l4+BVepHTpNJmbPy59TL47CfuuKmB6mCzzH2E
tjBAOHFOWao1G4TEozu3YkvYjo3zlkmlCPwz5KNza/+0uaqYkHcblH46aBg5DJGOB3i/QgtIL2NW
yLOAhcm/fHrmec576vNAlrksfjK8DmaA4k4AWKWIfhXLMTwV6u4MVzIs4JomdRYoVCuWiUTB3oay
ghCmJuQ+ao43n3ZgsZQ/EHzOT+0Z3NZnUAO7OAkp9QE7TNvVAK9wrbUsYr2ELZUMwk5rA4lRU9F7
dyB78qhx19KyqI9/9ERpu1LhB9gEuuX/sb1irH5mYto3S0Cb1efmPyOgjVgYgo38z3mR1XQAsMWu
O22RJEsFqEXYBoR9XkRWdWaiacEEOmTG704s4MEk1M1GjuzhELSnyJzecqiuAoffOhUWvueMLVLH
oDRGuoyWtNa0gPwTksFCJcOSJ3SRPlkvHMYfXc4BzhLee/ZI7p5sqfp3um65tNP7NoPNL8yjtLzU
i+ra9MFxHXbTmxDcT1OIz1K6dGsHsfrg7h5xTOamn5yUBfvRmQXKHGNK52z/1N6cDnqwN3eVxbl/
E4CFJaZoS0ue2t65kC0JKoXV+nLNl33vgy0A+S7lLRtOw2dCepVVLPynnOGF1bZ9Giw7dIyRt3eh
SPDO3meeMEvm68AJ+rh21myga0fpoTtNZY5MgcnGWIEkkqJCKFprPM0QdeG+Z+/bSc+oc9wBN4Aa
DtlQAmTCTtKLBbz3e9jXobVv6/e1HJY7ylN6oCX4JLdk8+vIlO0d+t72k+Q95BUMfvWYMVbSGGT0
lpCT7FU0xHLxyoFlO7gtPGcKxDHVqK2Ebn1iFJFHPDwm45aoZXBCQlKk+ONoa1ej2ntjM9cpIcPl
x9jYqrkMggpvb7wGGDQMNW3ZzBRsT0iDKbU+5AKHpY03jZmYyIekSQMaBzuQoTPr4OcxL3+nOq0O
cgXGYSpB5JyGxhUr1jstmKugZ/TUaW9apgA+zwotTAcpuHkpEHzSo+0h0yoAO+5smL1ZTc2CO6uW
2aUb+ijRIJN58dUUQbL8ine59s4lOecq/UZhHyjjMr7QF4dIBRHEu8ShjRnCDteGqTIudELFEb/a
FRHh4xnGlVzIkyr06oTFzWolDzQ8YQ9J2qwePTG67zlDbRtFAkG3YU8wiIZ8ctLAGWFMv8AhPRbv
psSYfD19SImypZAB+lg6wKxn8uL80RwuWSt6LzuCcL3kKaAwAWj28VjLv4XNbtHacqyixY6BLr8R
PhrnykoyuB3gvjYplgBMioLcDxSoJczFj9pd7SbSgG3rmyvS8T5VxjNiV7OKHjkkwPRi0QY1WB8f
NN7olrwISmU2kkShn3R6HLxBRQ+9paBz1FrrlocMmjcDt62b+nM81HMd1ZcuqYHe2PE9PweWohDE
A02m1hjBm93E79ebY3OXVnOyCbv2D0ZVRw6jXAGG3e/Rk65bozvWc/4ASwM7GWKNXD6t+TD6vTmI
/+jI34e5WlVkiVqCOc9hSW5Pw0Ld9K9Wnv4ARHE+KUmtago+RIvxNc9XuXpPSyYJvTt0YWgY63Rf
1rfRo8iE1peZ1BpuA69tuaEAAjgeulscE2j8Rufvb9NhT7iyOZywjroMhoy0CDW9LJEZgS+7eWOT
35gqOem3F62Ncjfa+WaJxhzI9vmnGYzdhiGH3UZx8mHDj79RmWpvPgRrgWkdYFFaB1ktpw3LebKR
hZ0ODx6H7EOQkCx6JXao7J3U3YUsglvkOkcoi2W4CLuYyT+ldvFrNhIqnMblkE7Z9ZfsD1HH3cTv
ZzVWof4ZRCIkEUIKX3N+AylJhFOFppsQwNW30BEhJeLkedlHZL74gw1+JJJi80xdoqqYdHLe3nt5
Hj168tZX/nU+BrqERYOO9orocRcUcwTPjk5etyHTiAY3oJb0uNd+Ald/QrPmy0L4S94gv5f+4Cgr
ZN6s3+k7PLGoYwfabLaFc5Odw7r1cFUZhEuDyUBfZoGTUIg4HTg4zVJFvGJ7DG0n8voBlK+CfXf2
Oa9rxhrF6BMXhi4YkRTmThTpd7eIPgQcf6kKAqnhheXQzZu18JqB/e+yPhJGRDSN+pz5dmsNQsEE
6xjpUjWWAi6z4ENujxqHYNSOn07QxsNWelBvv3gqiLp5is99zXFSbKbx1QNle+bIGuUFUqhTLdB9
sd2uB3vv8FKaO4i9iGRNteCPhbJ0HYY78OAfjLWAaH6ch8VuGJVynDwi3xBJG7kQJX+yQ+uyL/Rx
VBc3ONFYQUF61Emh5d5GIc8lmj+g09V6bsGXQwvy9SRHU4PzgrKNxv2STI8e2R6FUl0wXfkpLk6c
0RsW1YLIwkGLocoYXCdAgVyUtRNBGPNI+Sxt8y/CIAyktX3eWz57XTUSQpz5GG1stRYZq0Q/S8HD
LbRcwuwn6LK2zQjI31pymf6+OWcHXRCIchneV/ZvhMc/jE7UyQOViOp8xFtmV8mAfqSnZti0gXFV
sVI5sW/kwS3VB9wFPR86n2Yaeec/odnxoh4jaitexvvGaTEhf5CIzWsqh0WMtSmKgvWUi2N+K/P2
ZeAKgEhVXtRA/nS4RhXQ4bfi0Z0Ki4MPAnOZVudNyKLlBSwBryI25zgQU4nSmNcetjHf+xuwKYe0
W04opQozj5w5eD/Kx9FprQV2u4QNyyQaWSM/ns0WxpZ0SDV05dyh3ZfD3iT39HjesJyot8nq8k4t
sNzlWk3xdC9c/RFVoeB8JzuVIJAU9K36YTKqgT0jSWti0vbyOvVs7m5ZPYYtu/9kDsiGKunrAli+
DdSyONkfhKGBFQwxGanJfkfcgmNSzDIyK3I6PAzXkq/hfrHiAiij3A+Q+LkizqbMnL8aGf2N4R2T
ZWAwsMdiGsZ+Z6ahmc0HH+3376pq4gCdiwF5873IZfZvVLzVXslUs5pMljtWlzV3q1EXWX4SaGO4
IZhjRCEtJ9I++f5l5HQtGGiFcoRPVCprLXL515EAOIMUDIS7xDQzgnfasREwb/KbFuy8kHntgd3h
2kNNwKcBlVZGH+DPr8HDRjQa7o6Nlo1X+HDpK/MUFHmw574Ap/1qILoPtQcu0qodrrgiuEaYkkto
N87HdhdkeStkRUJbjld/kPC+iwUS5TCj4YGaxQve9G0qrlLqvaxt88kPERHzcVBJfuNHTgCvhusM
WHwq8xzXMNskWqr1XntSXn+9dHK/K8Tb0cTz9u7aiiaB7sfsaDTL9bdAsQzBVFR4CjzFPjSmFFC1
JwE+r7AzyO2wVPZhrQbcYLWtfXMOXZ8w10AJTPQAurJmBhDJznivo15GoZ3Co2uNENV5Rwf2oulx
1tS3SqNmFdkpj3kMipAB+SjUbLatLpt3fyKyj47/hc25SJylETtP2LYaBv4gJbGAdH0fW090d6bW
UDwiZKBf3qNs+RG0hr3Mw9+2G5bf4mKL81857PWEgMTPb9qRjPQJwU0fOYJBBNBuWlFnqTdA4XZE
iQbcUiBOSUhdPIa2oQWZhvqPiKiJtWcZlykka7kcZQng23EE9Fadlk9sNV73Mg2RjHigSkaelHWV
uSB4/+UeNKqOMInVZ/Lk54sKBSy9vvH80BedeEXABof6ML9qpYmH2d0gcdt8sMk2gP9G80qnnQYQ
jLvoOgxBjdu0ZlV/Wmkt1W2b4gv+F4P5FxO/qEBswZhDHKEf+VVwuvzmJmKUx2nHtAzKU5YgDWll
9lU2eq1OVVkS8NGICMtk/lEPUrV4OZWwAGOFcbwUXfwAOBgsCG/l4x1aHojB8ACiu7rsYrG5OTlX
WldHWmmmI6NqHbyi0Yw4X3ok59snQWuyOl8jbHyxk+s4uTSOgMimV9/T11blV2JccH+f98L3EMh0
aYhOzGM0q1/IDC4wjmJmo2GWNZPw9/SMch0ZAdR4jmyUIg8qI2UtV8bIrY39W+TgNojmwRcE/Inh
eM2lildYpLDf4bRFk81AU8QcottH5ROiToptOv3etzezz7jUYc5MZZTgY0TVTMn1SeZUX4rUush3
fH2NmT0/8wnd+T/3iN0EBwZQwh5U4CeWuADDlGTHrRiZMiNGCAWrcX8arJ7fnWwvyoo9ijBO9xin
GwjcEtmaHDYFC3Rdvw9nIoRXPzYeDOLZEiFku1dRnfDkQgO+kaP1oud6uOBu8/T+zEPAzMrPnmbX
dhVxw/kU1olScyy/AfucUGcEZdw7rQSNCgZXRzyGICwkGOJdZw6JXoJvmEhSXmkDP7No1XSP/qLm
nNHFZhn0RLK/bmqI0JVOp6x1L4PgWlhDnIqu5Nkz0E3j6JQWn6QrvQxQmxsqjnBd8EAaDqpQcdr5
1JHMYQaPBe/BAD/hvyeiZCsuO6ace4tcajWGnPX9kvQUsoW32sUHTRQbxBbUMiunUx6l/BltC2q3
bk8+F+D9hSosguRPwHVfFQ1nTfC8NQbEA0t9PCknKQEcARLnf9L3WGm24m01V1nd0pJIZHDA1TL7
WbfVoqjjRWaer0b4sS5ayBdyHmxp77hNXAW+Y1O6pTZWz3pWz4dTIBfpuH48gjhtwlkByDdYljt5
j40A1qxWRGYokmgzq3t/Z75mrJ2olXOO0bc82ONY184Zl+eoEk9oY6pEl0I5if/pn3mI+wl5Atsg
WZZjWCSV4LgUVn35GIiyXpoSZPQjIqDIWQUz9wUTe7rEdI3xj2UjF1QiQsRSfyRBxL2MQcYcOxOE
nFoql4sggS/RZf9ahuzwi4E7cetFNBPXDRzOCHzwhAMWLeXjc5MTtfrdsUjj8jq9Z9RXi+n35vu0
XdHTcN2mrLrNaTlldOD9db3TjOjPjjtEvzTEsZrprDUU05+vDuI3M18b8X81yY8dbImA1UiDNWMJ
zl3fH5FDbOdfRUKTaH3ofxX9tBpeJ26rTQ50JaLE1T9uo8dYlU1k5m595l1x6xETvCZ4sJszpmxR
GA9U1up5snkCA6L/CiJQdME9N1TIzFh4lKECF+CfSFtLPF89iOZQ6pNI22HRBxJhIpc4CJYyOFcW
sDTM8ks0qP3vn90u67uH8Mlapa//BMXjE5KQfVI+vsofV26GtQhWHYBLgpdlqd8hvcIhzZZoGMXC
JiLtgcUjnVldbbMPzbUUHRpxfWLIF+72iWeWqEUXwjTWIbMPvMvpg1v6li7T8CwmUBnyyTkrpCqP
D6v4dkZoAyfcXKJSxxZqlzLK5KrafQI8Tsm27mIxURt0ZuB2wrPwS9n3rdvP2kapOqTZRfFB4RWI
cAutHVYGrkkU5457eaD8VLz8aGLMihB3Ep+n/mNW3Q0hMeSUDBlVxJy31Y0qXpbUi6sjUQi2NFBR
6oKI7qTCJSDc/hHbdXvPIWt6tHHstAR9VlqYWL/ej9cA5xsSNCWYskCThkGj4jEnqzv4LrFKZsDf
UmuzwQu7F5hHc4cHWXviNRAZoeEaSzqmxnbqH+C/AupB4pOFIbSTykkfgLNACQxDUS1b3ashlkRW
HXf8yzSotsle+jGyE5FYVK50n2PojySnAHDgV+6t5LD5dGvL0QnB7yijf6aSh2uYzdM8ZQALISeq
9no27KIfAE/NdSgCPEI9wQYyO+HyoI+U3o6AxBy1YvPBPxbRvatMDbnDMvb2gX405x1UlHh779dO
WJ6YQm7rdg6zLcdePKsHBLRFprF0Y53OKfA2sxViiaUDPhnZV2Pms4jJyr5kAJslfk4sLooulekZ
ogx9vjcE/WjxdsdxwEcnnAUn0j52DcJxAxpzkOQRj63pZ2Apvn4JsbRTCNzYqo3MlnSElIpc+ENz
OI7enSaUMuARHLmbrn7XXsVekqAhM0b9ePvApxyS7sS8mbeln9zex7eFVne+5KQ1irn22K4Z0cT0
4QXnfYc8Zp0Rub4EsqMUr63RI/f7bl8in/oGoXwU0cS1uSPYuRlDRP6bFUNJypKSLgfxa7KU9lsR
XDHD6An9/M9ju9UEh1GIhE4/dq/1UTDNgTatVmthUcYgceSWS9PSuqsix88E9kEA0aOcnC2s6JMU
V5XCyBq4wIBNRJ0SMr9EXW2NyC1iuvmf0C4l9lo386JyK3wnwQBK3LxhUf51v5p3zlw+LPOYhRnz
nCptAaJP55UN4FSqWoVYFXdoLA+NQOhZP1JEJTKn44wrUVnn6Y4EdF1FYkm2Vl48DXwpfCNh4Myz
Zj/s3nG/QEa2hdkxQHpOaWumHTXyX0pBIcq8CbmvHmjzO0h5BIZ6szlpPMaVo1XIPbM3KC1kTyHx
jmd7bNP/gxuR3mrbR3rnFhvoUFyaUlDXCRKgR5dxdIVqrzvXRSg1W2Mj+kd3D+bn6NSRZFvvPiAr
tnkf70et7fxrtdlpGuWUuL/bqKNS+WTiz1mbGzFiGMZ8/VM4GJ3paLB53Ny/dUgGnwTqfc+yZmVq
ibpWqcjsDGRnM/s9DMGaPVBEhU88UJ35T1fYRF9sAwzJgDEDpzp6ZDwhPSB1bH4fX2t0h5dbQR78
6p+15t49aZ4GVVcgFSN4BUS+j5XRUY6GD+dHAS2s4hfFxox6rHyA0KVfO20Bh3ELjBR5aHCENX97
ZNlISwM0Z5N8R+SA3bFC89Wgq1zll+x8/J2jiAPCBXS3dGX5rZO5SQbM02K+lfqbkG34gvLbGjJf
xkZBNvphZXY+97K3+LP53jjHcvowYPwZXvZg0QRl68h6PBIgXF9fNyAfvdZQkVplO9iE+S2EJeXd
IpnE1Wd+P6mK5BmkpIvNAZoU910GNrOIIg26cOAV693gVDDu2TT+AKbTv+WffRFUjrRZ6pYovYgd
ItFxXe7uHTK1vh7KAS2H3VdPunAzWxo4PfPuT5dipuGIEgaHSwXdPfmWe573uv5rfIbsc2w7J51A
Rkd2yOBcLXjA+D3dSlqgRL+vdjk7DGGjhbzTRSQluG4OMA53WY6crgDKZFH05oWxY2R0Bwb2hyZ1
PrPTPpZhzzZCsPTWutd0zOsxTPoPKSl77AUYQP9XijvAibie/xvY2wYEQ43NSGLG99RDKl3R7yBD
e+pBaA+6qFqzTRFOeNPZGcRByUaoa4P+z58x7ltNmPVb7Ors/AF0R+qe6c87EcnAc68yoFIpIV+E
SLg6Hhd6TB1nAeyvu7lJgKh4x3UqQhBEIlJc0fXZQIsAvG1itMzHI/6MJ6DwgE2jiBGoCvHHaTCJ
s8ijI6fkBINNlhrSJkW5NClICfFSxmXNWDGHsPEJ+G/4W+cxQBco1lTabL7wyMT5zI8+24D+lnzX
/q9IHLtY2CJ46UM47EmB6KcBiQWy6iUAtEorlzfpv4mzLFepT8l7oGFgz0UxwW+Ok17UBCHOg9Bf
PBYNFjbl4D7h8f9Y6jq7PFwgyLExp+HsE5aXTX471wIky8COgnYbFYa/7mj6/H0I1PEgrEyB9q+Z
luMgwx10aJHOFx9CjjSm/HgdNOjI1IevIo7D/wSygPa3UF5s36tGeFVxLGwlq3smnncbS0pOpv1t
h9y7fkHsUE9jyOaId69+oBY7MFIHcMAV9xydgvvK+0QCNDphrmTfSbDGNUfkPAlA6x1mEW4z4Q2E
NC4aly1UKb/RNLm2NqugKIqXYtPzaF2qLxlZCyCGAS4E/LvHJGCe6o41G9AWIg5x9I+TIU5Odpp2
WMSFqEeL65QPvPKqwe84CoI6ZehpbVSsv4eECfVRxmPAWWcjVajEx8zMemyBlrVaOlOEr6LEn+k6
pLla//+ZN5mopH6uG0On7S+HCN+sA+LasJ8qNMhC3RGqu2t+mRxSSql664UWYeQAYz5O+eXqg9vd
fbEZ6huDUDD412XUKBxl9wn9Hqax5oiV9e/R6j11N3usXvjOV4gOnLkTB2E68/TF8eNiM1C5JaPP
AbHJTFmCyKDsIXL1iULNcuc6ikhw9XOCs7zZ3P13E9QSQk9nDD43ZAHDx/6sQtw/GgfnLbM+YL+j
pfywYnyO60PtfBLEG4GtvvbSJxMtq9qFfNwIR5YDdZHeXkFOLaWiW2028waujA97sckQr4joozKg
cAxZeV3jxatu/67cMNFmanI7h3wxuzrtskMHbfZbYEFCDR0EfO8UjW1qAZUQ6wbr9eGDRfgcLfB7
VMtd39BpQAcenfikrrvvDdznjffcei6pgSoye4pVEIgZTPOF1+HLgffUHeI2rcizUe/p7n3DGqlp
cNZdeup9DQxVDzbXUJhnMP+Zc/EICiaPifAo5WHLgQu8u8+HcaFOgh8zECBTTUGLqyrJ9xMnMHIi
KsVo4prtLgcdZznnSKGCbQD1QASFq2lbzwreZIpLFbxtOLSs0gfqIacKahnFjzJ4nBFWarAZIWdK
Uq2SQveJ0kLW/QNE+A9c6J+qjWPIyjxs2HCAyJaydnisgPFsVa9w47lzAa3WLdGNZIsBGZBPGn1S
TBSVqtN+MiTOik7ARLDVK/Wv8MekV2YiU7XBGI0bZgheqkSQVegHFFYfEMf1sJrKfdY1I6rEiaGf
vBJJ16Z7txrM2+dZFL0F7HCjrkt5P1Sl79fQqT7DzV/QV9jWcSR1olGjiQ5A77ZkA183qCgG/pyY
MTePUQtyMTWnOqyHtbnum9Il3K3vXiPM0z4vk55bWCNCw01+ziJDlIFB9zOfzJKToh4Vc4dCD4X/
1v3i+xbOx5T/rUSOPJKlBUXNrPfx3QU7m+nWQAkv1z+j7uqylz+APO1GYqt8T+Pz2Xzzwoarv9LZ
Etop4dnTOzXMdX7W2noM32D1MpwXy4Ly9VMfPy9R9fi3wxayhq4+MlknDIOKqTWoq4ZmDGJQ78is
c6nNbF6YVb3HRWy13Gib+n0QiznBS3TxZWT6LYMj+7UfIo27fvJK+LAhqvV/SgeS7ztgmzvunrMy
+XAr4z6/zSCGEIViFRNZHq1vqcazYFyW57SFQtFbOuOchL+La1+g3XsJ5I9snIhM8uT+AikPw3MK
tNqGnADjnX1hg7oy2bDTFgQfP9cYyoeSjHcEZvYTxrqm1LtvammmzyKlNMnaScBIdKbOgtofYWFx
RmT6Fa/qWzRy8g+9LXUqJBqGk/0xeg0kq5mtJBIy+wJoNtv44aANQt+dRkp25xa/WLuaMVTB84tu
dKsYo+9Som42RzmxO+8Nu7cWJlw4YDHRO+1wFLY0lhCT09gXK6Ijzugps085SXXRvAKGIrDDa12E
fMupc1ydIRzdhB/nJroOkWSLdJQi4RY/auIHFElzN2vDxUKfV37Ub/fKqLi+3kqRvvND/GlyJp8q
WwWljMCK7ELPUNHH8vT8OJVvacZk/IKCz/M2HOmDuYFOFuGSem31SMmjksmpI3QAfqtnupl60z8L
r0Ij/joXBWNzwwLFIHLB6IO7fQKV5/zsUgCIwjpPIykX1w+b0ge0Rvqv2iERDP9kzTZnjeZtm6M9
T+qRQzdnvl8GcVssJHmPnh6HEC6fU6AgzBt1OtZK82ssVREWOuu80uKmWlqcOu2LzHlthXWEZsaD
BsB3Tu4yGujGwGr2nZJshaeJrJw4qyBe7iJvMMDyDxWMqTIeofnWZ03m2FN37YtjnoGn0H7LBH7w
4SiJAlCr54i5GXmxI5scBxkQRydkKNVRneSctnb5OFI7/RpU2k9pZDW/2oALuSR/qphuUCPuEcU0
wAp1MrtKc3piVzX2VikofJw2MXU64DYWRazlj6NE3QNmXr6JzUWLwXsKR0PMEgnwCFSWJDNoPSm+
ws6sJH6gahShnTAF5FOVaLVmi8jTs/G7yrAszHLZPT68V1nT8UNm5wjzIkcG3uU9MxriXV4OcXlu
4auDHow39F2x8QW7DFWXk8qW+ApWlwmlToXRJHkZOnnxmrjbl6e1bchP6asYxc1TwV30NX2jnUuH
2ty2CrRgAXvz+qVd/kCnzLc4O4kwQGrNO4fa1/+1XbQpwoZ8wUmwsVdy42UrR/OAXj89tXHZA8F+
133AvSG7BZr1ebbBxLL6bb3zMIY1tUelrnVs5UA/VTKpqGOB6WmokOCXcxO6u1XySqeyB/yUXNJm
tEF4Sd9GemhiD5gTa9iY8UNluC1MvWxRPsBUm5esi8v7VF3K5HBKBnOVfIfDngptEiM3FB9PSYRa
N1UgdnK8asV/vP1Ddl1lPOLjSCK+806DP0yeb72Hzef6dzVsjuKMYUECHFWnkf/2cELwB1c16/8W
G1/VpnGVA5BIlvcz8k69bjtKZTECq6RHHtv7Nj5Z+YDPCDZlsFo/0fyfuZ7PxopcOIqj3eQP4A8g
BjyIPvaFXBpDL2NbQFu/pp+jTaf5U+8eXlIxOd4/SRNIgoPb96CxZlcQFtDi5uC5yzoEWSkiceDZ
fn4sJzQizJGxi6OXDDhq8kp8pwuwO2r7QiWUvOzsF7KiSk1qhxSeKEc3tA+jeRLcu8MOrQJjDtQD
V84nsMRkqq5Bge/IdlFuFoFxiFo2rzuIgIN2iYoLkDKxyZBRWZZhzDb0Fz44eueOMQnJqzG5Abp7
kFZ+zwxgX2I4wVt1FsE3Wrc6UStvZ94C1HCrpRSnLSD0K4AajdDkfAaMLEgCOk0Uvtohql5U0KJW
OBOlB2Srav7OG7cBcBs5E2sc62oULvuXF7y2hCltzu2L69OfRqCfHgTL/cMv/hbpAvZfX+LesA7D
ObYDngsa+/P7EPfBES8WUBQBSx2fOl3Hqrtefro4LyBVEhGsj9hK1qUuI9uyAxD635bapqfzDCYD
z5Ikfmi/64hZ3cGWFKoSCZQQ0B5Vj1uvcDzMLeJSWs/QjFrceFuFOwp9EE2TjUGUBvXd0PtbbFil
UZJlQDlkQ96SMm6A0ItjxqFuIX6qSrsCedIPUecT24zVzN7+YgPgHGTtGxBG+G3LYhhW2bk3t6pk
sx1P00XcE/I0utBRXgonEyzKoWUX+voEWdOi+MOBo0RrjIXO3C7RIe/TndpPfjMx9BbVWvRce2z3
s2UpreM0acfHgMeuNBZIhmrF57DnWR6CEX+eMguMk0eyY6x2fm7V0wgo4d3p4JGpQ2bs7t9XdHfx
TNLFqHjHYxYWj5PGgGqvqHl3tEw0Rqvq77+J7Ktr0M2Jr7GPNuVR8FjGiIp9BrLeoRw+XyhWvpTz
e6VR/3uanEon8jaspU5r4zLzfGdcPM1AqqjFvht+HtxhWCU+QmCKP8+rtPWE78y8EbibqEisYFef
bY2eJ+R0WS8suTYZy8WFc/veS5sN8ZYMzBSLIHLsJIFbSa1l+uBdwB1nJjmxNRdDt/OjK42tLZvI
EOutG4WHSIk+9LAwhHlazOsi3dtORB/aV6tOfnVR/TV6wUV7plpuKEPILE7L34kqdSzHfQomyYTI
hp7GLs08Dv+RODNAbVhnNzJLaGRHBSklZocccpoM9/b6nx+vW80yhsSI4yOBqzAmS0wAQyNgJhTE
L2J4egvSwiiVjHPam4d8N140RuGWo6cf0Xx/gztFFDasMLtbTXQ7yQ/8zIzNRZp9SmoKzAKHuMCL
6MBuwZ5bC2Hn76FhwwQz+sc9e7DyXvCx6mYV0Fv/9zLI8rebl4oQ8s/oSnZbgwn8wVv8HJKrqbyy
yvFc4xjZCBUulBRAsKt04BVgMtNAjXrRWzTH35qkx4DT9aeKNQy3GHh+mFdN69JrMEEz3ieRRUhy
ODab+PW2pJ8ciSDXcYoEUQixARFJPpAq+FDWhYUKUjNqm6DoLgiLYt9HLW9sPEsOSzM9n0WDZbAL
gwnDHMY3qCcDwJPly/P5ZX9oHoIkBYN34eWAvFJIWA8xspNEjJ0vfWBloejOwimKwM9T6f7JS7MP
rgU9dimxJHilAJzDPOhj53UBSoMZANZzLxyXHP3uUpIOz+nVlgdidaMOPI5jm43hZpe1dM8LX1z9
ouRix5ncXWqEjpsyRrWK8LuQawsz+0BQmxPANJpJ/MMTdY6e6eV1VjQfQCuSoP4joU6frF4LV0Fx
ijzxnOCHzp68HLzSdZDp45NW0I8dnwV2AqV1uA1OrX3Qgg9P3xJx0EVooH85rZCOsKpyWg1fxErT
P5StVQFZWjOFE61shkvpFAwzmn5y8+XIn8n1BXswMMoeXGfJcAvg4e7yCt/z0g+LmqHT8cEoHjWY
GRvAphyrKHoYt/Bom5wWZKTW58rXnYqzh/JOSSNoTNFPzLSD4XCiKQ8V23F+cJX1dKlOr9/Du/87
ICZotz9+OF50KvgzWYcBpLqBVehOLW9Rt2KyJYdV8o/xq3JmG3DDDjuLsefUHWD2dGnRk9tNFz3l
I3Fh7cE+1Tsg/vODQwq6/WhuOuGlAg6lelmc6N5pZkBK71uFFOLqk77vCuivhGwUUXgJN/KoFDxD
ecWLNve0NeqhVhwr7LdQpS9idmbwAvE22qEyDfgUmDJOPh7nA4IsdScvw6KLrHyEkrn4XIWCebY9
XakKNaVJ0Vxby/8Ku3U2AW9qzKdOA6hc2RkknT+zwnUrSA5024kIGms8wvmj1bxiVM0kqOqKXeaF
HyUMq5pNlxfmt9C6F5bGh6UDxyAaoActryZbLEARcTxYqTGPu64asbfdT0D859PKKsH34TJEcNPT
Gj4Tubjkj87umv79wJnWfNuftFfyZ2uh2o7bd4HCoEvxYVUqNMjpcRXSp1ucCQHF0Jf7ybU9KFB0
RkpN/EPm59z50Sc2NGZMXgRzPnvVh9iSa5f8r0n+Jnk1Zf9qQ1ruYNk7s/KzhDR9t1HAhH92UmMk
KQ4AS8aRk1S3rT4OxB2y5FUZJ0P7dXYkavi5qJCIflDC5v2GPgE62iEemMfV7BYfIaXMv0L1Mrtb
e356pWh235xwfn0qPjPTY/J/QH/EDJbVA8rq417AofdqPJODwMHWYWUyQgb3IdngEApoLUWhfic0
bNUYMsheat/0zVFOH8pjiybmh0erI0sY2M07u2qhl9TooPS6rgCQ37VM1WICNKGuu6OKCVMD0Rjj
qCF7o6I8A6H1DecC0lwhyusRT5PAKQjkmznsT7xYJlOpPO/aIHdA/eX+b2UY5FKVyYj5RbtTzJ0c
CPz+x2cZLSyGFhaKXB1NzSCj8B+bBvB89P+cxUWDLrvgKYMek2au+h5CF/e4FW18Qb4LCuaKYVvt
F4ORH2Y543YvzNGVDrgbbuZvPzbUV/KDZjfY6UFMdopvan8j6ekk6cofGhGI8asuHGgVjmqyay3H
cuUi+uAvzNqrRllpsJLSzLTV7uxchn4lF0GDjG5AV/r+kZ/XbW73oloIKn1C/d0EPzBg8m2ZgdfQ
zLqWBSXn5b4kDTHNFFhwi8YLZ+WxFGWU9cWIHQMo0Hkr+DuaxWNa9zwR18UuDLcEgBptPcHac9uY
AJwD7hNdh5x4mLzOz2T9MK7k0IPCUwNMFkULg+4rHC0Q/7XqQ9NSaDA6pUD11Nn3fz4kxyD/epKT
RJoE0zdhng33CF9f304PPTRQ2zl1357Vwswv1YzTKhtVjUANqiRyLx2CaBx3yyL+d7o32ecwByxR
N9o3hIap/f1TizF8hxKrnF5grmmQR4PfAtOrKQk7TkpFU319+5AfNwOCC5S8l1MJ8fK8HhfUt32B
7Z7rKNCRJf5Hafg3rxfuP+cBsSYytbmfwjb2nxJ1bYBWcWUHOgLu0Q1EldkxTegt9obj8QGw4uH/
EHh4WylUSYk4J0QBYn9J7vA6w33otfBL4eVAye3aPrgmj5yfwoYP1BAcq8nvVQOMBqFFT14hKTQg
ZmPFpFRfSOJWbibptEsSYY2+llo9UrkPQjp+WCLI2Cs4HH+XrU6vQNNWZQCMyFXQjf2ZxsT+OCDz
6EjvHkO4opBqh7kAgCWCPQcSECig0MlLgGTkxo7HVorwZYmkw4KFerAF2gaAWhEOLKTV+WJmf4oh
/B//iWBgV4kawYxXi2L0HQZ0yN26YPx9zWodWQ2nJ5EwCKpax8oBQvOwhQLTDuujoq2mDf4wEhea
Fi8cVRno5Pv9StPEyFPs0Qs3rANf3yNY2DtqDSXz0k2QymvYqWvslgpRt0EiqrCt/0MHBHYM8wrK
E6mZREn1xOI/jYwLY4ii2R94ruwU52p9bFyQMQaK5t8pJvbcYYhfq9if5n9fH3EeV4B/gX0LEgo7
XJACnyrzATPn1q1Qqw8aOHr7B4/sRIVIZMR/3xjLPECgbyhBd+eOTSfQcEiY3XQ/GPQPm7otNBjM
IBFUS8tev9q8WuMbsvh1HdpoC7yBh1KdaL0Ptu6YvE5SWF4w0XtXOr6HOw4FYe7gWidhNdHgebAG
94zsaAegvuFshhar74zOxkIepzea6F3fZSevTkYepfEAC5ikkqGOoZpEbph904bhicvmDM7XNOEL
L17Py300xEf615i0WQtoJhsb/dad74Z4aR0MCp+q3qC574RFyyBPHfJzlotnHB03R/SOfx9WfVCk
vbLmrNlvRJBjKw8qdoUFIaqbH75GWs5CUyYGRafeCXeoGK6I1VW4pIWtwRD9XivD8lcCCeinCFBi
vnkBbD+iimCp7q08PC77XLR1vfO5plk3sac7AzhI122bPf+RY7/+dLC2BxJdoluelZINJU7YkbCb
lDFgwTmiZbAZ6X9cerpYwUq3Te/CZRj7ZeAFsPtujLscskeTdNBJEi37hyg/V8GV5kc+7FUwgH11
yAOjkn1tBz62+YfMvWSsvhIOgG3+8WrBvJVPumnacMb0Z/RediDljkWE7FHUOXhCMfQkBYG4FgyW
H0CXh2IVZllHzR+GQzDN/sN4ukTnQ17TwIc1Yv9LadQ+hh5rTXglrDtOzN0Crg0teasxv5x1i8CO
XDTYj7o1Q2Df7TjIFhxAGVngVHLa4GVnRNasUz+VFZs023FDcT5nHzddEuw7n2YBUV9p7EDRaEBR
ich3hQSnNpCeTN7HqJvsCbE7WJ8GOHO4YTaCFICF83xTM8i8W1jGAeaqbc39yuqE0gexbw02Rbga
u+SkxC8KkjxiBY1NMQ0RwthELWeV0xEZsDSZBXTllKR9R2waotJ6lp39BwsmVk2nYGPh6tXldFvR
+FbPPHIrzL3xW0LYqH6vClEVnE7yCARk46tmf/2LvRG2+FmMTs7wd0n+nXLffkSXNf20ZF4BFuJL
GG9J3I+0Aov6SNHg0Qjf+Tgy+UipS+EI9pqOjcerSY4YyDMyuZkhbpgxJiKbLyjP1smCfW1aP3/F
vlqOCOi7jsPQRdVLg7Llz7Td3G0jmcj8iOgTRvjR1ZjQHxmotYh4tePeZtV4PRXnBWMB+cKW9pwf
v7ip3YqMRvVumDGv3OXw+EQ+NUvc4pnjMs0XgQr8OvqClIdmN9+cKKjQogXxfb1CGfuenPJ1P4g5
S/SE1uUJMK0XemqMRqDdVgXhEqvfGcPOoj4CJZ4cG6uJ98UovurPKcX3IOgFvBPZeQKUM4nXLGKw
qQ2vX/l1u6qyinllb16Tu/QwDSpyEZE/xXMOMIJK1hJMbFbqFcsd8gCSWhCBuJgRVe3ye6otl4N0
BlZcgFh+aFGbKVMMpKDax3INaRudt9Hs5wNcbSPAZN26wieNj8CBY7Sc1RamwqSc6gmFZVDuP0rq
0zSVDnL2umkYiHZDvwNhOqlqKUNWb7mMXozWWjXE7u7wKhMn5VBRq8EBzbC4pDxoAbAezGr/ZUqd
m6CIOoOespzZH6PgiLvmj6XtVSsDsC5JzX4dHqsYm/fTFiqpRS31oksRoynYIv0AKpqS2SHoFoOW
diJExe3fs/IInjoaHUeN3ZQeVNSljZLUVgWnkq9FNrFSsREEwe3qs5IHKDmvjmOHcJyQhrR2FsO1
GmKQskAmIGCw0TqXvgEryayWtyf+lr+ksQ37UbMqtovm7jTFD6yxdnBir9DkR+1TmjyxWhnmjBbI
vHoEwKduLQYkerp0CYPIj8NmBccaBb5oU66Bo5beMlR71zgzoyodR3roGXUmYIgQHXn+PzwY1zmn
kFx8CoIWnE79lN9+Jy1MPUvXwTeKgVRd7TcKemAn0Ln3UQsSqeRI10So02SdRgFjN0vUX2/CQMRS
tbduyJ3+7i+cY90LvTK/1iuSJb07+URhRuij+D4NZXl4t2H09zUqPRnV1t7VwUwELSs2qBO2SHjA
81TnZAW6eOPMvFL5DAqGVGjcrOKvJX2QNxpSirUnCiicCYIbHSr9IuoQhxrUjr+3WswTaAkffSd/
Xjf0pVzm4et/RAHqYvC6qt8gpRSO1fFbp6LdOymcpNQNauSszi2+dgGSnlvp58+rfTxaY6Bmm7wC
8cSjK9sMb6tv+NB+pEGU+PO6dmTe8lQKQ9DKCev0pZVRisZX3jRjmN6FEB8P2Fj20d3lZ2aWe67I
NvoXN6nJvnjTFbRlwAUGh0YLyv3Z7Zrqry1xeNBHK4M7780vLauMkU9iI+Hyq6JaEaahw4VbUggz
iQT6eHx1o4bwe96aGbD35ByAaveC9/C+KP0m0BTiPxNo19UBW4joKyqtdXtlCEXrxLSLLIl/uQ/w
4YVg0mjjibykSHkPT/9CqjUyRWNtsJTi2yXFFnKlrP2WSlSA+DCWfeKbdH3PrBY0zqcYTNT0tPoY
rgqfEendTjoLNop4R4y/ja57xb21HpRwqTLjs+tYBbG194LVnuZUS4/zSu3JJtDI9z8VVQqVd6r9
v3c2PJfXoxTYcSbWWbTFazpreGwPTiBadfw/OzUE/TCyf7qcOZxvWjOqDx83ez1aBLrf7s+zzlfi
D68HxklLWDJJwzLnas0Ba2TbHhkV1fsVMdG/dtbYGML2qXvF3H2aDszY4WOlTO3CyQyfHeb0VpR+
zLWf2Ur98Y3RLgmdhcX9XUPkbDE91v0KUFYRLlZQ94vNV+E74h2KhcNuI1zfSteXzCuqeo7N7ML5
ijxS/QTpRcQYjTxSjwkjg11DXr1Xiu8J771cgeFEjdxAWvATPkmtfEsh27vc/1vpSJAq2I/fu8gG
tgEKxd0vnUXVdIRX0Je+ENlBt8UkrQmdElLSixNcwhjUwCWSS7TsMJg7A8UKtbepwHQFePhvrJ4h
lkwwZywkmo+dD7dguCYUhssaZn1eqFFi/CH4ozj1EgeuTxxQCaDW57LRJP+zzRmB8Yt0OPS6POA2
COesJLE0WuXF1KcBijPawn+6zmaYQJf9Wl/Coj8AzOp4WCrttYQXgnJyV/xD6AxDFgOap/WJWqOd
9Ueq3UHazYcGEC7JsbigK9Eg10HZCnh3o1azRykekmSCIQOx49Y02F7VJS4qcpYcQkYkf/SbfM74
4ZnRNesnvxSpvsso2X0n3vlyRg81nDv4wQIeh+ziq2NDGjJVfYlZEg0jPAHf8eRmu7blT9VHSzdV
9XOd5bh//yfuq98rQruPvvHILQKTl4E8MNk1EPP5Tiz/ncPqnjf1zqzHpjgV+yQhwpIjbZ2CcjTz
fHkJVsIVx2e/iad4Pus3n5CL92l52ad+mP22d3+fom7t5+u2cIrDSDQoeVcDFWRPyTgSOKE6zVal
z20MrD7Ucct2U7EKMLQ7n6BBn0Mb4oveIWCl6iphkVTTa/iV8UMEDPuv1biLQo8KEIF1NMB2AbNR
BQv0lXtvQXWyOzVIH6Yk2TqspWhfaZEcaKurZbJ6N/U8ihT1ZAsMCq+tq3afw/OIo0GBiHDj4pS8
8GhZGt4W8F5/NlMTkn35zEVGGIS3Pq/gCWQG7JY2ENlF0kEGIZ6tUxvOk94i/Z2dUejOoKFCxOiV
WUnyYcMJOX08pxxaZxepJNX3kA0H+8J/PwH+ReHy3oz8W+scijlXdbDqNcZxqsbz1AC6f+LAZLm3
8UkuUZYeTshxoLPYA4XuITAvXBw1ECYSeTcfIp0SqJWVIHXbxsyqXeCc/722ENqrI2brDR91Yi9L
cXC80iKWDxG3KzPKuZtwL3VQsSC2NjBZACDvbF7IFmBRKQgoNJFjoLURlziCKm0oQsN2UDaG0PrL
nYJoP8zSF4IbDd+iWpM3hEt4J1TO0BenNjhjynjl5woEXQEc2xQMQAGFTmIAHGBd1abxhzCVsDwx
/qFzASe3JvswshkgtKN9B3VG8eZa7rzInZPeWGo2sIfb+uX7hcLQjBDSJ9kRkFEAwj18WO7g/8WR
fGSUk41nT2wepGiUCie1M8+oF+h31qekengzksRPLiDQr+QNVaaKbnUC3dNEXdaFYby80gtuuIYo
F6W7L88MI5EPtz79APPaRyBfEftu2f9aafCjdJQs8biPYKvIlTSkd67WlyoYiHTv45TXrBW55aAB
sxLl0XkWsV7mpqzosQF2fkFuXCcP29wPQ/tQP6YvOVL2ag7Ovr+g3161u9jGcWOK3ek2erfwXNSu
L0IQqOos62G/7CSY6rzObDLatuhAm9RGwaGi3g/Ves9oQNz+5buerzJj7Vy0Dge0Ncv2wsUBFZEJ
IFuwoV0oYpX/ZKRblx9eAw7s6kBvPDaXPPwTdpdUeGUGkGT4oPjWqPf7MaBlsNFklYF42GjOQ6Ic
z0jCMLFuaA0DIO949nwaJ4ZbA/6lvA8FrUYwuvaqnYuHtawpLTTmxRWG079EOrCutJuOwYB4MG4P
x62TQpZE48/xkxuuc++JxFj03fARPn8qLqjM7ZZVY6TpbQf69hpWAfGjeiXOj+yT4e7lz8/DWb0M
CJn3k3Srzcka67km0RDw82fOBRG+BFx650ggwwJSCeGDRGODPDV3aMPW+7Vj0IXeVAPB8emJ+qez
6Cee027eZgKB9H3eU77l5p248DuyhmKHY44yHjzE0AYGyjAAmjQjcvB8E5A2mG1WWb6zQNXX2uQo
ozSocNNvCdxVgGEXq1JxdjIM9kadBMaTjDKwadbICBL2QZM9iYR6aURGVCT2zh7sbTW2CYF/P+M5
pB/EapyUUX8gi+WXOfvc2Rrzbxc5Cp9UpZqG8LX6alorAW7PihGWDc0hXNrjtGJs5NB/RBYcsy4c
GMXyiOYwSbR7VxMu3N37qm5Y+vP8F/DYPRAnALISsSQWIsSUMZBbXvCi1yHSWrBx9HjVSU0c5D25
sqe7sAUUgVw69cLZsDygocoaDrFNd53erauBLb+lSowJDNJbU/Wv7brH3D/28urVALFQ9FDhLdTq
XpQ0Uyu9KGMLS9qOLAPOU7ySNUCryhJLUi1lBBYgtZJHP1Oxz9GqfSnXFAXT0pSwfkwiE3atWu2L
2SkHClswdTiWnp0Wo2xzefbXWhAX8qu7QhRKFzeneOAFvJvdSTsVrXHYXCP9BW318LAPKVs0DA0F
XtwgW6ZhnP6mruEs6Be5vAWYqSVvujPSgPCPB3/2d2d3LsKb434vmlhmu8o5TKqv82kJC5+TjBoe
6H2WuZX3NRqWyhjKGAzcHriOJjFRnjwtqZGiz8sfrjchfdo/tc1pPfrbyWfsuPXqLV6Mq/6dGrF/
03QKHmxRh7qycj6o7SvcpYRkQKopCwRs9Zwp35mZL/GApjJ9cLKgKDOvzvI9pU9XhHrxOpmrr87F
dQSGcdYa47JcHZi+2/d2dEnSqmi3S9S8JyhMbC1UZLkWwkaxnOltuEbLJ2AcQwmi09YsdxLBsQbK
KtsI9DKHhtRBR5pjWGGeuoYzfxQvpF359p95B1k39VVGFy09B/YEn7VSiR3+L9BNEpLuUo/mStmp
0OxHMaxgI7s6nrzVfrSp6+aw55JNWOuX8NEz2bvun9VwTGw2v45GLhCntn4BIig2S6vZzWoLFI8a
DfwqhguC+OnKCaNl9LQbGi9l2FG5bH7UB+KMYW4FMG2zoLvwy++h19Qc/cbwZOE+XOut5qe39HEK
6zmWxHARjTZ7kwz6GYAq0+ZavgFEYmkOi2QHjJcSuHFk7GUG4Rzz6sk5DTeNTtDKDxNPlrGJBbfA
CiVYTP1BeNr2VrLy1k8aePlMsuB+0CNPo1v5C791Kn3qG8Ur4D9MrAeVIdxLgGsy2TBmmin7D0Db
FQXiGTfcmRr4ufaCSUIXjek5pVPjB6whOikZ55IehB8vH8wIv2JHibEZBbZTBiNW7deHvVFerzvI
hBrPheLRN/AblYbfti3w/b2TAI7iOIME0+Nky2m4fgnbgAtO7T4WuijB+WQYg5YOluI0/jM+SC8X
ND1PtT466g+BW3QK9JBmm4hq5irB0W1NS1c1h2mYAjkJzD7aBRboQkZZmgWULPTkscQ/bTZs7Dqe
8NzyGiREXNF07NXx0m1t6N1nPANLlOuHL81dmAH5fMvKEasDlzOvBsI6t4BeK5q+uptdgZMSXwIg
thRaHmX4y1nEZ5v9I0bl6Rzq2syYf5sNDl7cRVY6zsIXuQj9KNI0V7ifeDawoHFMtUe5IWkEgMbc
GosOdsBvcTw1b+XJxt4a0AnRMT78VtPxf9XztGQx4uSrFTPUHIgNXtdux6qy96BfmDm7DWEtVYbD
dGHmlOmKRLRCGbJSQhronZXgtOH+ccBOu7JQaXUkMb07g3J+zdNumNgalReMWv5IEIEdIPmZp40B
U5/ZKcZPLUov7ZJbYz/+lyC1YVN6VA7ILdoOQlzNYhAZi9PKcoLaJgaZC1+ze3bArCCPya4DuKg0
Dt57GBNSySOkqIuTadjpSHoAqbnOzJ6wQOeRQ98Sbzm3KV/xGJ+BUkrMcLUC2zAMlT0Z6+iERkZC
a11V543LPYCSMgld4NrVVnbLF473IjSFPej+qk7X5ggdnfWPGWxdgPkqCQ+sg+Amf9uEUmj0XX0f
8LxWpQpv5VENepLJPOINiwURzwO7EwBXmA1mQ5YG59BergQEPvwiamXQoJVa+ZO3PVEtCr5Nv+/i
j0Rwrg35/vMcG3zfGrBBHGxvIRMHsW4Pj443sfQzK0kbynRT7VIxz+yht+wOd1QGlo2XjyjpChVl
FL3NLAoFJV9BNZdjk5VuKkHeZm84Id0HQtokJ/DOGN+2Y5M2NxWwu6reg42f0TkTHvdI2l+L2H+q
mnKVsWoVUkWZXUhSFFyhhvkmWJkllB6hvnbUymImruh7W8ff8WGKGKolaVaB7WyK6KErDO8wCqQY
UpSW24ZaZrwu8fLP1kQS1Hq3rWr4C6ep1w161Pe5oNGbub1P3aM/Bb7GDiLywZDnHNM9eLDjfk6C
iShbHR/VFr3WlcZByiifyFKS7x0ad78b/sGUL1EbmkZPDdO5SmEgVMyFVpcqY4jlZV6ZFGvsQrZS
vn7SyL1bHH+R6o6v4Jra+V+rJa7KTXuQF8aVYB00GqXcN5MsQjKPQ5JpQNslY+A+nhu0cTDB5IaV
PAo22a5swHdACE8Wp1+74q6AONprEsYqhQdWLeTN8UaBrgrGsyuG9UJt/2qc3/dV1JeYjw+p4PVm
c99PMbSC20slPaZDnjo25ix4sjLgiqc/HLFM5pmTSR8qvPYXCweBykOllG5ajVBdaHZUUVwbNXrO
uFhPs0OxB5ANcYmwxMfU/M41vDXuJ42rqY0nLtdaiRl1XCAKbeQPND6LOHFoNthELF4SlhK1qfq7
rOL3DgKEImFEdf4n1sYhe9lOEAubfhTLI2Q6bZH27QZeRdtxxQr7RqJMSpXsMOjBZ2vx5Y8ETNTF
YzeC+Sp7zX5a70XwNdaHGXPFUlmokZDeaBRhCv0UwAQ65ln9NJQGIILZjN4WhTz/Bm52GX0nqtUg
MWwtY3dTX0QsvkZtyBYP81C6GFmXJ3QdDrHgtzcfDBapm/sT/701I3Csw25b+fKmpxlpwhSb4uOE
Hh2yTSzvPedar073FP1a0pOdq7qQeOhI1U+9DklfLc7JKgh7lxCGFaIoZTDU1eQd9fOSwv78dgM6
SbrRWjJrF+j3oIj6YZ7hWhspgmZpYdjZePCm4ok+HXeg9EHSwrEjaDJ3nKYa+dPV2KxREDfUD9Yv
0yaFUuA1CJpnCavlWAb9cHjYZ7ct9I6Pjb45OFjYWm55u+U3HtJS5KBcD68q1L5jHBBJNnKT9uLI
vr3Rqt7V3zQCGLv6NkC1bIlGfgflC2d9vMaCnda5COoSfbKR3LzAnsaDO547AYFSQCaT0+nyBP/9
/jCTeYUjtO2qy+7JdDgzqZj6aF2v87Yu0+zMfQ/YjxnvgH8AMBWhUgRfPWzCLKS0PUGdvt9knqZE
R1zukszpZt75yHTR/Kjy4hHtzb7e9DTBrRl7W4GogYxrSdwmbpwCmM3tDcQqUcPH0fVBiVCHKD0f
Dm7BFrWCIAjLrIL+Cx+w0t2p4BtiFmHBVLTotcXtKoMFnRInRcEIa6BpkgApb5t2PQHhOVfMOp9X
LrTEUqZUe3m7owD9wh84lA8uV971APVzmu57GI34FPg6q9/I+Ae7QOpALR3ZQzYZVcSPF4yJkaCI
P9ef2ElUpB9e9ssIA6bQPRDxAZrPF9+8HVjyKmv4nC53YKb2TveV4hSXFZz2pdq/dQ8bFT2egbfY
1pqTKcwHo4E23BlvGXLUSSFUa4ulCWCareWGNtMWrwSuAcOZysw4wjOfUWHr3noE67jFbQf2Sfbd
y+UTKLZxO8p14oYccRroyGNOppiObVYYeKhKw2R3jSYcPR5M7vBbhoBiROLSB7KwxXEpsMrEAjqG
jBIMoIpi3v/lWfkreA9hS2qOtE/JwV6twQEV7K9BDxcSTQOQLLvvTHt0o+2I2SkIsBZ6NIEMXMs5
GUtcFnZ4kfnOGU6gs7R0NAplU0orTcTPjr8cYEDhoDC1NRmO9rdXGgQwoe7vKDCkCkGRgv5UWdFp
Y3rALvCGMP6tpp+RudmACnQwzXZ7ITdiJpxKgWxEx6B3mNdgEfmdNhYJtHy2gizzLeOnJ2eba6Af
7Q2msbM0spCW3SjQjz/5epw6hmOUboOvsjoIITTA3e/SaQPqGAm7pnMSESLoNR7JUBeFCEs3f1x/
KP8A6txtSI2HpTg/h7HIOIwwbi2cS5weX3kTAPZ0zs1caX3txYmuQFvDUS2UVeTPVS9oOaaCf3HC
zBCpsgfzxUW9NaROD38eodgy7cimdnvVZkG10oeExIin5ESIzT/7j2QLR5CEb8s25UG+d/KUlMdZ
cGo5zhbwyxKMe2fUCdQqhPIJNmX9smMq643RdGEYDqWmnc2dBoQe82AX/Q0gth0d0EZ3m2M79+QN
p29Pf1lP97V8ec8SyKdBCAmuGdDYv8Q+quZkv5TzEZQuty0cFgTN/FX9RMKGrpwtB5bx9XlMt1EN
/hRKyXSUjEMw3a+C8GR5DSUTn2NsKzLji+2jYVDIVe5LfXpwXBZy7hfew58CgUyzo5+zcrtOSnCY
FdZIXYuK+1Q4T4NbeWIOd7vBwK7uOCuFwMu3FPIwmhGRkdQok1qjubKvOW9+Uej3EQfaWkI9anJ8
uPbNjZ1XJqpSOUD72lwG4ddplpUlmCYhAZ84QCIqzPQKmr5W5GkdkpW6XcKGZ3bJMxotnCspXK+Q
koVoL/yM/bO45lGRPWWvBBE4GR5+TYMndIlOkNO+9mx60cym9mMcF79r3aNnXz6cyuJ+6DFGuiTb
7VESPLkiEhL0KB3niorCJeZDma5YdVGlkr44WOUusc02vKaQMqTpeL0/MC0yWjpHr+kk+cRXDvkx
F/gB0nPdVbBmXbG2G9IA/jdOWOpkNmrsdzr2xvWmbnhzbkoUthMNmiYUUuzHPyiy3JJ8xrjVYzg9
bsiDlTldWXnI4HmLeDCOYmhENM+tw/TaXU64F7mrcgHNYe8p/Iaj6cIx2YZQwbuJ4OsqivIWKFEo
9gKkJFEllk9I4tYLS3F4YwdFype84jPZv4nZp3ZsSdtYJlk0xULfU5BiO72poR1H2EpRr6bNYKxC
m5bM9DHhlF5oldVCCaJxOtIfrMYGA+bDpaOZv/Itp71SJpA1ak056NMZZyX5f9CYkgOFkdCSO5Zf
18leI0as9v6FVJZldlyIazu2R8BgfG3TPRqnGfQ3uzxKwmSKg1I/CBuvOU+jl2kvNQbJYSPn55m6
O4mPTLmIad+ZND60uG6npd6BaN8RQ//leHNj9cKEMXEcVaZzlnbLpSu+cylugCkXPqRrTiUfQlXQ
m6lli+d5s2sMNKrMpNI/pq68xitD0GeJ8ZpCRiYeSyVtVV0cxIXNQhlfnN65AMcvpJSf4T0OczBR
gbBEraavu1Udwq2zwHtpbg2ii1/0iXxb7WCCosBhGDhVl0lJYmFOlPLj5OnfqUoEk26TD+JRVCeZ
G1SOYrHLCvYTwjrobVobNEiku2fzIrETvVd06KhdAfvK7XiZRbg82FyddMVDrNbK7hDj/A5PRVBC
jxh9WOKK3UsE6M+IDMzGo6AmCSp8X8Y0hzK3PV4QCdR7J/XSzSjZPOZLgFZPSgbK8ZiDW9fMtFDd
xdoTeyeILZTLFyWC/dOXiFpo+Fl6X8FdOu3YJIQqoIIa0YIj4JkuNUVK9P1WyZGH/ePC70kX+vwd
iy26KbRndTMR0perJDBJB/FK1GNTCka2iTBAMmDxrXxdnkeTJ/5bsXoVri/YQcG+yRT9yjwQlOuR
5hYxvex3Uf0Otv6ihyozXKYq73Miyf0bDo9F5sruxb12s3yC+VxMAC7y6V2QCg5GnXtvL2X2UNHX
rs/1N72iy/hKujMtorqGpRNCLZB5/7aM9Or1mnMZd7unoVkvLC1iLZXEd6rXzxPX6q14G6nahVkj
9VzIrG2AS+Tymba8z5UO6fvy4bY/KyLqibiRE+7FKFgHo9RMT0o5P8A56ZtprDU1gtrKRBInEZDj
Uiy6HrQeSv18nBnBXA9RZ3e9mysvmpk6W1xk8qKLzwG4q8JV0fuklElK5BCsi4jiHKz2PkFO/+3K
//uJ7s8Qcegy5dvtWRqSaWKfg69zpcC8j60bPcPWRI6xH5h8RAj40ew+JMoHXDQjLl5ZAsEoCkvZ
Nf6NBQbLa9rOVIaDdoawTKS0hA2ycQHAeIJ1+Ex7GqfVEvCL+panMStOqvJeSm9lJ9VLmuff5acv
LRWE1lg8q7GSwUq3bx9KXjAXKTe4zybiXNImiz8Yc5efGTknmP4gJ6j+VZqSHM5oLh8H6J1Zzokl
vsGkoS/wDlX1rrUQQzxG+XyidKIOb4mVAa7ep/HYuFHWUNLOWCh4+Jmdy+W6tsDwRP2y5BJvGZpM
0OmGEwtMw3QuAAKV4pCrEUkhrXN4k24ITwic7yDAbnOktrrnnZluxrer9fc1AK48vJJQ7ahpoban
xllbKXka82bzJQIiE3z2lTitga/E8gP/RjCpJAvTZfRyVdsyChJEA+YEkPYrGe2fyXbKcI42GWD0
lPV1Up7Y9T/d9kpSHW0X7xfL/uBAIE6bdEByzbJ6jZoSDmv6ZhDe0KQt0sP68GpoYZmudnl9nN99
iZCQnXJE0Px64gGYlBKm1zBvBApV4v9QohNVKfIR3IIgdUrhZBqO7+wkWGKvIvR7TPicV4wyCEHJ
jrrmu5V9vjQxRCjA2QAmUdWefuwe5mRL8zVPsmJF8oH31xX2mYcg9Xo8MOJLRMH3vjsSeiZBv281
B6rREvu/umBQglkbLz9/bUIQhRURuXqW9xBp79bJd6gQnCJd8TNA2e1A10Poi1Nyc6cm2DG3q7hf
bTqMSGsXnSQyBxex2G0Y2jN8jxOfYC57X/gmkNT8Krb0O4+a1BtaNBw3qzRgYMgJUmDykly2E2g+
76c9NL56JHUQrCqFJOOPWHBWPocJOOXS/5vW6Rundv4WZqW2VUgEZxH6ZHrQ3wOHb+IVN1DzoTK0
DM/YRuH5A41S+hps3ziWYwSZdMBYzd2/sY/99bfBfJfkXLioYXbgKh4xD/CN2/1clOoKjnMtSTYz
QGGXMnZbAANXmkEZDM4fw0yNylzX1ZHiufIOv/dP5Qz1RLa9YVZZoMhFKu+LfNvAVEQbbpM2JgTv
4xJWr85ImKCTEeXzY6qolWXirKQPaVnug2jn/5bu4WGjSp0WdXwkJVSlBTNfM2l13AtFzQshDHg9
A7hIDZowwzUsHyRr5pq6MiwZwIymv1cJnSsemkTZl/IPiy9fzUnQWxe2RRviodEMerlGXdiwFQPQ
cQZ+pRQ7yF07XPC+oK3t065wBgafdAOPMZb5Y5yuSzNjjffKFt7RKdSOhTxbtORDAdQcX27w9r04
KXJh5aDkZ2XeYQMdQ+HBEnIQXR78NgKCiVtyDTkBKOfqfhZeh0/T8OlHf/veBinTpPwh6X98pPW5
1VckSRnhT2OmaTHxaguBraKN4KTx21xyNMbDI4M+TnJ2jzCTmpNbwH61kq1YoEx4fO6zJoOhVJFT
qCoKEChyjXj+S0ved5OTvv1TAlChjU5MhDzGKSAaZv7JyrRy/ejYigrXNWYLFOQDA8YKjXZBkZf1
H818PkicgYEJfPWUryDqDgVSfonxX3WBaPJfb7Lb9kVk8HeVDhF2590X5784Tfiqc2EglsG2M+ur
J2tL+T9Bg3IZsiKZE6LnmibABI1Nj0L4QUTm9/LA9SFaocz8DKnP02P2j3bpOv+n2f6IiXQfk/mW
rFgukrquZqG34K2+lXUdOatbHhNtIRQ4GRXHnXbA86VKaprYPADQoBi8YtmFcLwMmZJtLKY5Mj7q
oNRPlHvI7Rph59GJ5FIeJ184sotPwMj77lFL61FZHNV4C6dBvrEGDBNlvvqYv0HOQ1EllmtpvH3N
Sn4OhPtFJF+wKQIP81Y4i8TSgkyummzCwG+I/Z8dAMjYtSFK4CL75eyUWkQOqnrryQuroN3emEoN
YVVkE3BgVbc1yxvXZ/wQjqMqBvSdE+Ec2llFrnJYuNqu94dh0ztPtSH5b7DOXJuL51iKKPvKVekT
ye0BclZQaAb14ayn1THHcSd8iCXOBIaGH5x6/X5uacNKeyMFjKdG+PCTy1xsFyA+oQzUoLN+RMSp
wDUZBVixH2budF/9JvhsI7/xd7Ch43C6oy3TGw4SsPdN/WOEvvLzp2dst6Ei6OHiXizMqbygQRoG
U40LPsFu3uJ+r+sCZh4UY4aJpTrRqyf3dOXP2fhBoIxDZEq1DbuZVCywbzblf1Ipxoza04n/xdRc
AK1bzij5xTHItpLyZwuguzVU6h9Nun+EWrTHOwjcQTm8ZKKWPXn5hk2JM3RrHWfJOGxdZC/DWLIB
nJfOtqCo3Fylm3n6lQ7oe0ou01mKjRXs97wwefd3PskrUKXAe/uxZ0WB1Lu51H5zqHLEtZYQfazZ
dHC+ZdqSAYQXUwCQNn+YKTDnRoJj2RVLVBefkEAYo9YivmRerwKwlsCN42AuMWQK1JfCNOGYLkGj
rnwEox5/boAEscki5OZb7e4yuDm4hHJH38K9UEm0BAwl++r/RoriuRHwqH8BOdmG6ivCa1ouI2Cw
rDF/FBJXAemkO6ePEZkt7F9/oQr2wohHK7/cYDGu/qPPaO0KDunmIKF9ErVw4KDw39pVc2SaFTEe
a2gdeOOI+hnt8cJdzq+aYZ75V8sXWDNQhOnliKkZ5MJl3jJ4AzMf5ZLElDZycOfExBIn2YBCbWcy
OpYAU3OK7NnbE/s2ebV5cjkp2OS5RjDSEN8YNG9P5nXC+a6Ft1id/LxCMT+vFM87Rv2IEiUDYgMk
KH5+3Jk1twK7UsQU1S13RjKAe96w9YjPTJYCWUy73AhgC67WOfZ95tcSvLJoNTFWtCPNzlcdJ2SQ
0KGd6kV1/r/hSFz9qFnT/WjJNnRUnCls0j1Gs2NuoZ0Wn5zT/AfleHLLMyN1tXeMh/e8EslK/5Tu
wmhpZxbIQijpX5C6b4dB2ZXVrObAhnZiawFW/KTVRPvCt5esqYXDQbEcwQM3XcSxskCrPJJWxO7n
l2/iZavTzTlDMQZxxLPJbp9ptTBBJjvnPD2Jj1sA+qfuTDwqTFuchpEet5m7x/hJKl9eA+ePpgfT
JZXVKtb1Y4I6G2z50ZdaO8rnRkgctarcdo4AU1qYQK03IkuK0LjXOTKiyNPVjgHVNB3dy6uvBuBO
ym4yQFC6o0XdImLmS4ep5i9TljxTRqTlRaedr/8Clf8E94QzheQLt207hUXXzkECvY3BQdSRLhlb
oISCidqhNCSQ/CKvY1VZO1/Qf3GcPy1n/E0Uo/U79QBk8cpbmFaxQlPw+rSEOtAClqCIRRv/Mgxe
rln901r0zg1VP3KwAEBiLQETnNe1MWC6MdvQC2RqbsgeTY1L3M9QEDBe/z9oqDUZdlp2jw4/jw4q
/xdlVp+n+jqxhPDhnSpyHQGyycc25mSdXRLuMPEGgb5RIlTHzzdvCtFOeCxr81mv9YWoVkMTc0N6
EdvG1X32K/y6sJ/sx+FQGgw2/bsRlQVQ8TjRk5zdBxkEPyNj6TzEIF72lQw996NXP3LxsyLdhgNT
8MH+4Zd4DwVhuIAhtlG2T8vbJoUk5OVM/Ohev7n4n6fjOEdWCnWVQuuW8geK/iWmy2xus7DVXTnr
ytur7gjxOXcqYGOYBDnmdZAl7v8GWj/NzmoKNO/6kfSySSLeIHLWbKrhwvvGBupl3/eyrqdluM0/
3PrfEnBsTvbzl9pUEKLeoKd/8eIrSSy1OYxAjWskNFKVyhVz0imj96MRkYvywDI7+zb2lxZUoQPw
Oo5HCg3Kq4VmQIkIQmBtKI60WVCMO1iw/35y2oFrsXTAFqjRbK2xA7Rnv9cUSCjUReo2M6WC6xv1
mCnK7R/I70uMy2xO7ZZMwy0W2des8OAP1fRYzakmL7g67p3RvJPOWydV9ibiBVk3lpSV1RLQPKX1
UEpwiRmw0ZIZXTrJ3sdbJc41oU+h/cBIavUMOxKyz52MtFsJZEGLNhRJ9JjeIV8jaFnrlIraWuza
jwf5/LIf0RWJCtKsJ+lt2XtU61R4BPtf2snMCa5D6HLsiepVA7wCr2MV65z7/r8lwB2ZGtRy32d2
E9nwoApORsot2DPAAo2OjZ4ujnF2tG0aOT8YEGD/UpSgaE1Aw/aHt31HayQdi9oO4bG9tLLSdKEo
lc3lTef0Ba/VF88KJc9pbhR55yTN+cWqj0X+R/zied4UQBitwJ37orggMrvxQYNGhVQwIW3cXB9s
DXlCYZX0eqV1EaSk7DeQjnxRQIM3RzPjOmL30BoV6Ghijp+/4eYD+q+hWIhsTGjOzJIddh4jBca0
7GJp/qRZDOokTNlp8Pf+WfMldvd8zZKcQj0yglD1Fhn9FQh4Uc3OVYX7YjoC7mKW9GoQGpKiba+j
0BIIER7BFpM0MPV0k3U/zNzTZoyNrCdIA7xMBTQONAzxBHwbOsjPk3xVsdYVj8clie1vfBJrJQ4m
8pwsqrbbgizxLPl9cPRiynmvC+YS2I6nMxdR1TuDvMvZ4Q9ObnIxhMDfxJnbBnZFS/Uz4N8uq79w
7C+XHSLJdVfJFXozlsizG2hEppKpMbaiJqB4EXMLMx+KiIIbdZSMtcHk/dfuvdPN12/OSjK6XUJ9
zs4uMDE5r/N1vB7F9EAaE5pBfM2q3DC7eCvc1d5O/BorXgGLDRVOshkRytPd90T4CWJrVYgDP7xa
oC6O8EvZ/+TwtYs/DaMmhZQizSU+f9eobUs3JYbKS9xeCQNi/HALYhCfyOiRGnN72+4oQLd2RGuW
VtJ+wsQyakWh97P6gOuZHpaQXkr5l/FOdjD8WoIQQdkbm3Z1AiFbYMCFRfOWA6DLEXr91Cd67Q12
anpW1833myc2Wcn6FAYTL0D9NG0Ns9M64JF02GqrCsWvUpnNBU/FGohQy1PB4w/ZzqXWpZYQcTHD
pcvoJL2crqOY1jjj5Ro3TvDsF6jrujPS40EUsax5Eqllgo7zdx7qmbLBoimIP42+qXzBY9FiyWzh
xQcAgjoXNWMllm09innFUi36JRqKzA0olS2/GIk6UmwjPHHgEAISKOhDguclo3CI+5EpqxZrMFna
KgWivZVlrjI0yUJutA2kywK4TJrYjsyNymS9U60TQBq1iQ1dC10Xgx8Lsb4uOjg9wRFEX09IS+2q
7QHeYvoudA/oNX7fRzaGjm6X+Cg6vE9K9C4P8rVEHX/VOubFkULjIjsCLrHdrZ6v8X8UusD955kD
O97HUHpMeh6Vtg+cTqUVRg+nmrTpdk0JBUz7dkWfmSUypRrVAqmV8/jjerI3716EIRVWy1DEeYQo
7DIJycQkIybqoD87N5E2lDEPHZ7bTwRxO7Z1cOLOc21s1H0hTkzaPPaFAFpADzY4+uIvMpwxVw05
vQQfLEiFa6MidgUXqCGKyfFhAXD8PRol5eWDbP+sfsqWqgItBOC5sdIr20vycAAHRPT7QWlsEOCR
ezj5go6DGRqjLCxRkQXRcWPNRGkUi+5hyfdbQU1LqHFyC5Y6hyLuRmHd7UU11114rbH55wKv0YGT
fey1zFUyEfhdsrH+Q2Cxqzhid53QGnJvbrNbZqlPS3T00ipPeazbC2EvQjp9SIiV3qVjq1WLdwtI
TKuuhP1xbWwwQRENvqdxvV+r04bxXnwbrLolAsw/PfFWcZueBoE29p4CPDGzOTlbjDRoHuio3TJd
WRhq2ytj44i43M6TCmKcrHiiaK/X8EnywRGaXGbsX93bIKajI3klpHpSFP2pM/U8dL2CkedKyGx+
Rd/pfghC7z7ILV5wzSWDtm5aFuobvyz2K/hRISHy3UwHCivj3TUI34tqtTGxTo0ExQea9JBzsxZr
noC4WiDc7sRPoM6rjZDUQ+RLew5bZivAhq/SQ6fa2AU2HV4XbwqmH1MN0tizCw/J+YevAzfyMtmU
F8zs7+cYwS9EAphJa9nB3VZFy0JtvnupMyZzlztdgtjnmRKsLkjGdV5AfpSfakqxUioFm5lhEcv6
7Rjj38RFPWDnnhfbG4FgrXlgO29hThIHiZ3DtyygDzPWJ/48gZHAmvd82Nh0tjVU1UDRdK5J9iFS
Kv5aXWgP9Yo5wH06mMgg1n6Ww9UcZ5+cFz6qXA684zOH0E3V/h9UZQRHfjpaCdwFCdHAbL7m2WWg
u/xSS9mgvE4FZXwKx/aDna5G+JjilgUxuviGpEpeuJEWnIU1jIWLpTu0GVAutLAxnfTE8CayTVPU
bSQLVYUy5+lewZFmJbTwYrgMPbmdOkOW3pe1sxu5OHm9c3fwVbpDevZbwkQgxcM7TisLCux/ujh7
7BAZBMY7sARNmY158w619J+EpGShppjyZDqwXnkeD6VwlwtDHyOBRar4qQE2R89Kvd3jKLnOO9HO
YJPhDRtG7CcYOewmAPFmVmac9H4dctdHbHLYkzVmaWSL8bjquVxKQ1bjZxZRlO3AhCM4mOAaZT+Z
/IcX+16YQmhEJ0XrcXTI3FvvW3gG7SHbNLdUHyyMMsc9u/lh9rAlg87CLwOM3LBBmT9UkeJ5iN6f
j7GeFHvYKW/GsF8GcLS2RpSzU44m3n95zL31j9pAzwK3WkZxfh791UuThliZMuofv+cd4kjIuLu7
uR82drkd5+RZ0MR0+GSTAh6d1pY0nM2ahgeeof1pKCQrOTt14MMcFDXafSgjjiEh7c/+CFrONiYU
LTY+ot2Is1KRqar+93T4S10iJ+ECE3BEKS64r0p9W/1+DCBDqYlDU+7Le82P9+9b+fmQJhkUOdDm
PYr5zrp2XwthQL1BNzXSQ2FVEcRiLXOyRWRDn+8PGQiS+AkznKEfFM9/k3QtibYcLXIilVyNmhtl
l/Gb6VKsNVhaR+BwGaICV5FRpYI18j27vGQCygy5+rAxWGI2BRT/GiXrHg9bA2QQRNe5X335/LBr
a5GJI1IV1BHDnqjEse0zkZBKxMQybeCNcOS8euYHiRk8VUv+mlz+1/WQhmng2AeFrp2l1jaIHtBk
kAST2aS9K34E8PVUXVeHSoVf4JzcDoy0oj0ATLACj7AYaxnvfR4sxXJlSQ2zDr/v70eFjpT2UY8D
dxu573ufHxIeG1HBBT0KZ+CHr0gn9ehxkv7aExZYrKgNY/DitrmPv3JPeDKhSYPqEG/MBusiyOE2
hRX1+eVXRyyiKIVMbto35TPg4nIteaBZ7GXvaeAXxNuQ/iYj5SNuDffcsB4XaIuozA+rXZbIIJ0x
J64h5fVTMaQjMTUzEdK/G8f7b9V6V9cZ9RpPFyQAGDdLDE9OSlIwEKrqPLhv7Q3asIXDCoS7ecpG
zEkhu7im4kQovHzi0u4TB99jZsLPDXqZE64j3L0CT0Btv/cvZx38ipmFOMl+qYLx5/ulfyHKz3Gn
DqS33um9rFEQ9GrMDZ3KMG2lbjkTQowwK3GfPkFhMsjyy5sHPeZhIpYqHdd/fqAjBQRSABz31Z7R
XkbqnD689kPmaj+MhRIVJRJqdumA8+ea+UbxfsZD4C459+Pf2DgxDKkeq5mUFrzlKyJSzRRfaHBt
BEu93sq/VDV1KT5fnXslUSryFF/Y/bkgjsnFWKEqaiKV83VEM9t8nfIGyQbxbrYXheKEsljo8Bnj
jKJWKNOGBwSJemzWNE/BJ2xNq6u6iUc9dIEvI20fd1q87D6KNlTPxqjCHVS84v+WOyizoXpPNCmW
hsyFgShvZoUtVaNDq0yAtaDsWK9VFVr5Bx9Et1iN1sdLebS+vTHuA+UoAWh7bGwovyAIYpV/4uTF
g38mwcYfSqs6MVxliGmK8Cu7qOApB7Zyl6RAqKP7mONqFLDbe3XWwdQPtw17lUaI/Z7AGlr+rjwu
lWkQ3VBO83nOaCNbQL6UwvNup3j5MHlOGGWRu91jqUAjkZSeRE3u55EB79L+BEl1pY5rUXOlpk7q
XqmsMzjyZMmVouukRyd7AQf/Hk0yTErEWw6vrnwaKcb7Oq9X4L2DKC4rU9ZXOz3PSGdVAUCIhV6E
1UHHV+RD1iiLsAfTBz+NySlF/+M4XeOyh/KYo9Z0BiFlLGEKgUewF2ndC69sIV1IYagJT/dcTSVO
cLp0TCy52RmhXLCA0fO+rEgAkUW1XAA4ZZRbEShNALFglbFOnjzgcKXA23hYklr7Af7/Zvhnxgbi
jsedzNqXC0mc1kBoSFjaO1Hignst8tP4IbWjjI93QyXDRitV9Ca/w17dedNebjooAgCxcp2rv1YC
qOC0oYIfHC2EWbL48AxTsYjprj/QeJj7LuP35OpatRSKmn5ohfIiO+wG1VFT7KJ5G+x5g4EbAyRr
RBS3gN/JwUJG3ql90WpmGoGtyHqo6VMAlueOYqwtQkJoPQPIUnvWsXvo3lnSFniRuNftvck1zgXk
coxJfMxFaT2PSlkvdZOE4U5GvORMqybXwnnc08EyNCKCu4tIfWuqx/VB/ZTLJrrsjwm+l77N36zr
8UemFihP6kZ/ni06isV/ETRa6hpjb64GSYd573hQgIKNYPP3NNjBmrbTNln8ltWhxAViTCA4wXsu
CA8IVdgY8vu0hN0rAFX+veiIbxKAXBDkzlbGjYAM0WTIkNqQ3Le6rIaZ4GUWmuAExsFw8Mq1TqtZ
8xct9d+nEcAI0lle2Ah1QRypV/T0ZvW4p02Unv5LmWtf+tMZygpiUFSjYdSyYnWgldV8mgvyALFN
dUykKgFlQKCNuzQMDbXBeBo9Y6fCGcS3ZDBx/IXRBEqtRugBoqZsQ82FWmQfVK7JDYCzsdlwePVA
yq0dlB53ExxhSXLEUv5kjvCjkSusTL8ynL+Y3qvap4BepZSc1LhhdVkPz0XzBZgYY/eoF9UAiCAp
+8UvqXcX0zcR3jd9xg4tbUvTZ+Ls4Hmo/Z/tWFYlh8BhW6qvJrn+UNsAXZJJtWPOhhpZqPIIHILK
npQRld9eYxcX0cso4iPWD4dS8tQhVBUKX/TupAIbppJzLAJe5Uasj3CFlC0QARG0OKga7UuWQPJv
SR9GJwvo8OOe4CjhBQCQKKZjesC/ZXsSad8VkH4oBs09SQkanKIT58hawcKsO2dhKVLoORByxDTq
7D+2rbtuNy8JQHGTG0GX4oXeWFIR+ZJ8A/fCh4ixv/I+fdnMtdLYQE3m9xn4IjGEUwYVgeLNtHrt
usdieA0VVowKiFNxlkNRKNCjKNZFqwa+z07XYCIIPVHCHAcCiOHYxKc6h6GoCtRwBUxeS5bvlggW
kljPqixSMFg9sw/5K5Lu3f3Y9FuGBV63Qa0+jLF7D41VkVi7K4KzBkhqc45fUIsZxgYSg5SNXrN1
/uURfpJ2C5Ma8fvnDou19HX8WecmeCrHp1NcqGaE5fw8DqDLJXGKSb90BK6ATETbAJOXxPUcFWI1
BjWQKmn/vbaxAuXNTTW35DfUQ9Ad3fosIOP+1vO5QNITerFx/Y786vf6qRk/KQbI4KJlzZGqLd5W
loSixdQSiI0exVtwCGSbaucgMu0pYAJLFbPmDUaUJxgjGM4l2R3GJMGpkUNpuUZvG4sPAxEw6Irb
chJE0Mk6+ewCbdmzHOKlGV8ySYFOyVYQisFhHCW4sSGr0zJQZdExAFe/bnexJ0qpoVlCtBhc//aP
LSFJKKJrSdIxGoa1aIxzjCdpixgeyHY3kisIWfa9hSKzGik2F+y7Pw+jIQTg7Q2hVJ6slR9H5+wh
x+oyZ2YzCEXpxBJcMV4oQbIHVsPveHv80pb5krvCiMRcI3ca92gpY/Yeiq+5jekMee2Spg8O7Z5h
R773uzSl/ztLn5QABsHvoovCfRI3z6bYlDOULGLRg/zcdPqHGmXQPRYfDHst/+DAlVdk57nT/GNX
VydKtY/6U/WxAfPijEphuszff/qB54HSsBpPoscMuf0cDrBCdCNCEJN6e740FSvsaMr1UPa7AhBP
52B9lpIyAWu2bER3Dgmjl93tsPRpT7cxe9lhm62hT7UzmXtK6CVck6pD8eQFZuMxompvIBECcpYS
SiytbZCC8Qh6HOxTKvw/tWZerTsK4eA41Iin/1qnO9jU/bUmAbSidu7N5AoTfvICMpfPqmIk4sam
8zORgNQLul3p/NUBe2FOoJx5+KcmRhGHKS1dB7f92wxKXhZ3e90sQttn4qtkPOglkh+M/lhTIP4l
EWhYrHkCHv+ArotiFXrA4fc//pw46hYAGrk8ZVoDCw+4s1wwifh9QUgbttY7xrd0r6sFfNkR4SyL
2pAMgcdSTX1UK7rrKNFBGY+60FfvWg9lltKWv8qbqGsRWtf7ENJZwenahYPmE5+9QLT3QzZ0b0OZ
Nj3H/V1xJAU4cX91zCy4iilCjAmfl2qaGxg0YPLB4B863UcaM7vELEB3VsLe1fOCYwAlWEE8cMLA
YtQRNlz3QRlIH7ozEnvq+RlUr8bQt9h1XrHxf5Ah/iNNuWS6N/ex534GsSZIAt1xpnOkYs7VLMjy
wWsdW8j/8dqTIrwJwv3XwW/3CqINfmgxRNo3o9u91L7PpJZ1AyDArJHALmfwXuZu0/ehXK4j1d+w
dozBPYSKA3dQhQrO8LPwY66iZvCL8/Gknr7QmknUJ03PSja8awzJ1RhpRcJAwF5go+d7W1P7DLBr
ry37Eerp6GRIgSPsDSeFtUnlPpub5tO7MqDPG+9r8XoFpe1hi2DBkSZ9vlboX1UtIyFkgxiV0Nqb
V0QBFm0GpJ3Je9OtOEvk2HK1oyb8JBJNwqlWTGykCl50MzfiZcLHsQOvJa2piP7eqxRszo79Kha1
kOvdsuFdlMAyppiTxrqD2sGBW06vIo4aoaUqO3wkSvn+aKxVoP+bnHCyps5MHx2bG72imFoDp0pM
FpJU6r+hDxFGma2LFYJ7ORWG99O/O/+lCkUcGOPd6kCoMUzoaPjK2YR+SDtXTNwQeq4A44NJ0A9k
opVdLFzix+t5Bcp9aN2zGKVPITSxCoqikFbNuHYXq1FJayLUFYNrLL/kXEstpNIOI5uZa/ELIzCN
HGD1dC5dRT7wYuro9t1NT4TUs6QD7U1aza1cRvK9xzon8Tvwx5miaFej6DtYp8bZiVW7rx0yLlrY
beBr3ObLdRkdcSdzz4/blrVa6C/qtwWJjMyO/RVOryh6qvOnYKkboG1/tAy2bae2NgQkQvcKIPKW
vQvYmFq8cTmdu6kdXbG3eGL+JGGUQJdyWtH0LZmq5MX2b1XsyzzOFXxcaLHYAPNbFM6UZLyVLxPp
CprExGJ2KSV0nMv6m6hVvw45VNMG4fUyR8ek+XEIBzbFMezex6U/HqeV0zh/TeUZzcUENu1LjWEP
J+LQ/WeQfgn1gVxCUd0wLwyDEE7xy4HVcFytgk9ZALscNpzJQwNFV3w/33EIak7CA4wPSLVSQkTv
cZHbg5IuvC5Ew05qaJdEb3KpJBbz+tS3/ZmRceTb9mS9Cmh1l3NcsA0QrD2HSWmKjsF0yBAyrUy3
UDuUxeSHw3EYBlJpZwDUipQ4ARw3ZrrETlsRocx8piiwqpWmRoRneoiwBMno6hz5lnj79gYkdBlt
1am9D4mlKLu2kj4Co/K2vguwWb29bwQhIcZ4e2RkKYpfIb/P0x1SY+pGnULwgcbFEU0XsrnV+6Ll
3Tfgh4up1HHa1M0s5IF6GVxc2dM92BGUdJqaL1eB2MS7hRWwmKw2FdMGra/zFLHL1RF9XgCWcK5c
bL+deMBL5vmzSWCiaU64K74jbj3a5E/2HdSVi/SalwOP7CqqQEpl+g/yxE49+EejD3xykt64NNMX
FWmGb+q5cD6sYyNyGNBs11i8GclIjJu28w7G6yqFQeQ2J7m1BL1+75shB1kSfSmtg864bkVBR8R5
clkSnRpvcHcxP2NaOgmY1h8VZpaFevG5pIV9oS/Ptj2eQ9GH3qUP2/3usmGHW25IXbto/WZIomlw
cRPhQsrMen3/CGgOI9qFO7AQFRnwJRP7570t3Cf5Nz+2Yab7IQSl1xoqLVdrGaucdhVohZRU20Q2
skgD0rvwo74xnFy+VVkrDO3YxcUKYsvgc8rv5raZwYSB5jpTUzkwxp7kT4W/ck6rP8SkxO0nFtDp
6ui2JGYGZs46InQGrj0TE+DQQcQnd0Q378LKVfkdpMdROclU5cJGy96n0wG2scTmNoVCCPF0pd+Y
E4+FoCRcSYfatleAsirzRZyl+U1j34YBYMnpiXMZ6qx9A/YX+kuModgo2Ltj/1DwMOPdW51WQHst
L7kL0LWmyeZsisAqR+kUIDlQAmficELKuTTJ1Zix0xxG4lxGBM6eMjSooB/zjBTI5EgutlG0ZsKb
mgZKd+xZzdjIZA3N/p4yxGO82tfENswYaUpYnlPxmH/HA6XUdLFiTrmEMXX+hIYUIlWpbxh21R7m
7t77II2uoQxGwjJLupAHEwzQCMXo4/skUY7Sg81G5HuRvlMYUOqJAcS/3/gdqtPqyvDDCnQncALA
9T4xvQeQhsj6sJgCoANxrqTZeMPqhUwqZM7BLzu5hvUEg63ASm+oj+cJANmLqxlyHhePr7Uh+RR0
a0BFk0YfB6NqNFN3/MgLfTVJeZSXNgK7euJZs6UGIIS4BMlaHM/lABMGgpzR9EpOaP9Wq/9LWRAs
hbFHrw3chOwF9at1ZnD87iQuUvt+GNYwBdVJ9ECj+fW8j1NNtjPSJb7GkoDRGGVnqeFITkBt2riZ
VhJNtBPqiOcjLsSGmFes1RJ0PG/3jRbfh8k9+kJkgjDYr3Yj0T+UZ9DNhqviW8ivquP9y1NNqud2
7Z52jhUEVdLhk6GaEH05EScZoxh8ExtoSxBep4tAO6fa5uPeejMmqpoPeRWLKawxmIa4J3WDO1kH
6GqQq9M1jsVHFxq96HLSn3K0ViBj1u4DQNQycNxzMAmbwU/AmxcSJK0nq3IXnxhYuWa62A4mfivM
XrytkF80iF/HYsXUiQQ35IiN1hgcyOFD1OYB0uy8jMEdN1AGbOiHdvYgQQZNn9oqIUyeEqmT4WHw
byC+TltQ8A/DRBzy8psMEqrYJztm8gJ5+e+ktyyUUhJIA8woeJ71jaaPxs5I1JilHOLRg9SdKpTT
eeThMYNolRQV+LoIjK4V+C3G2se3ODZMumAOVstA6HvVYmszsOILP0Eq5WmwkaxBh0g9VsnwFD3A
AnL2MM3uSgy9jSDrINeQvWtUlWSaIEyOVqfRYitPJJN3txRGA6+X+2u/sHt2sCMg1X+Xi6Q1s9w0
vhDFodMO2jHB22cNDj11uYHsk6lg/6Zw0/3Zp7HsGMGAPvZoeg0KeT7Z3af5Ec60KIkXojV7bys5
IHrOGr1vq1WjV77RzT/rYYkiF3u/37z3tsIgR5FjyhZF8rqNNcr+NebPZsaLewaZDt98Mci5OCGw
FiI+6NJLAkk5jBp+WXqs29pEnWd1QF0db9BNJu0j8tAMksffIfNC1rIJDwoUlFQnho0Fr+GUQszi
xELAe2QfUHv+aRZvnYTQ340fDlMw3GRXjZMkIkq+Ycpa7qS9Zw9ODvbPPCWpYpwj/pQno/88Ma4F
b0yVImfiWZ/Ysu3d0Rv4uP2T6I/eeX7Juh05zE89y7sIvYjcJ1QxBquLzQK1S6z3/tkCdE4hNkOK
kdJHvuygzrJUmWFS2M339wx1TPsajQrKNusPgACs1IBRWOzrFl6HnsP0S/v9971YZyCSegZm/bxT
6Ale475FtA7h6F+xkqB1vPQzNoB9mZu3oPu1bI8bfMimMU0FQ/Mt0/4YM0nUGBytb2d3DGaLS+bv
OYN0YgFJNbiPElKvOdkicknbxESpMJDPbE67dSd7+sMYb5I+qbX+Qn8w+cwdK+VueG6YS6zcKuDQ
LgvQwdXY4i/e9Gqn/Z68/ZpLV/wUTcpaagE9NSkVHXJRPBFMy9yLQ0sSnfHs0Ag8WkVIKqqWDZHq
RF9/IhcIRAayU/807/FfbFs+KskjkpSB8KSg9xUmIAIBrlIlyl05a7s/4f4UB7MuvUZTPaE7KinR
PZxakcdZTDoUAxeCF6J7ivMhSs1XHpdMqmBQ95ceMfXXwfwAMMq9Rs3eWl48VKRDcVr1VQWp7weR
8PM4Abwt4F39/0FWXmOm8b6tGyIEspIUN2d9Fg8cjb+aeliNc6V3f+Jmf0HqVMleVan8IUnZWkFQ
mD4qkoxYfpNfXyaesx/IMmtok32ZijGKmTyTLLR2subF+iricVNAGXIJBTgTuY8z7+N2jIQmFBof
901PDNAFg5sF2tyTMR+VesrSrDlBha8rzRi+A2S4cxU6UjWdTtjgnIWzCRhqoIBQiXan2IG9qrlC
WVyQa4Z9Y26I/0sNHClera7UqIe4Eq5DsHLCLdhlxL9yeGFM4jFeszXP7WnlhFGR/hpVhzltD3TI
7qythQ60fGZlfHgzeFQdARnz8YCTJVW+0w2g5Myho8lmqlZUeGpdW34XhHF7pXZ7FtDoQ635MVrE
anLwcElwrh3I7Ry3M99tkoae4wVH6PFHHqkM38UZApYwAigw+9VVJbf8Z4AbYv8DWsvqOdjPOATH
XyPLnukuxLAUooQxiw6G3riXII/ohg4t1dnI7DapmAFh9O47eoINvd6u02rT1ewelKxhvKfsdsIt
HUrzPaHKMT9+69qIxU/4RDSbpLa8KbYMP6RgLy5phvvVNnBPDtaAaOpuqy7t91OJLoNmeiz8UZM0
M5omZDchajtX/Z+V0scP+XA6d5roiSqM6fIQWKMKG+98WXPSpYh3Ql2n1DU5N71cRyfyEBhClCpL
zdktdl1aTs2N7ugsXpAm9a1hSyxG/VdqCpuWRuRBDXtj1LKFdKTPFEOLDlc49bxHIO1PGA9yKVhX
SIHugr5GQUrAyncasgJ9US17CQp++cL9/4Kfve3e3IuJFrOauDlQ0ZPhtFuUmiKZxX21HIyQek60
Sq3hRVWupBJfA0g0NPj2fzG4uV6yEn3omtmLpURi1Fsw1bEGeImJWMdJh7HrkFvh6ONFGZNI6fEK
BJt8Det7Zai8YCCZx8em1alNbg1oycTtBhLjgMzihCo98UImeXkWll+zFVv2mdflf45d2yjXQ/qb
gRS+SXg+Cmm+uCYoVXqGk0fGRKAVnWQJaYP0ogFX52+/T/XxvQPRMi7C+/8an5SUf4oJK4xoEg/k
iLw7r+cXLw2snG1qQ1UNuz8oyCQwaDhvujNu4+8OM8DCYQ9UzDXZ/56MXOuSYWqZ+YUMkm9RoeRa
EqSoVtBkbFEwOn0rxCL8GX26bOIRddv8n5lO2aKaAPDxH2w21yhoVqyX5495zfi8sKQt4g6kwzi2
t1npOHNq86MoVbSiddGWjIvJL2M+cHj738sfrUtK8/V6PmpQCStXNELf56ejEStr+PR++V8CVktS
90sVEojNmD2td7snYfpTi+O0s+YcnU0vS2KEaNWWgY6OyNt/KSkpvUoVuD3dlSuW8UX/OiyyPg77
gjCihfe/z6+VHdOM8uiFOHc+SDecRisrPw9QSF8o5/gTZIw/ngkhsiL+ODQUMOYmHKk0QiKG0HQI
hgMocunEaRpQAqdqctW4S0P/HnWIvEagt6S5STuZDzokso71tOZjCb2AiDaD8lSSzUuE8xsuGBHC
6yx+DbeaA9C7hHlGnwhvK+u0bW6woAwZ8s/THNIjCW1vFajIxhktZPSt7jcNcfYCoJyE/9e2TpPH
mbh6upkGkbLRQhVle4dKW3D7CmeAds2vwGw87ZjyN/IZvmnQKp671/OWvve9iIq8N+/CdPnLL9ax
p5TjaE7nlFAytOzrOm5EjDDRpf6EL7lZ2OsGFkSZf+O+Jdq5nvPL+SPiYoGnqRcOZ5zFDhxR0GvE
ZXjOqcWpPItUuUnVf7JGjw9NOhiomM7YthEir7p6M59ceWe1ZZrplHjPugSJZu6vXKYwFAmpYLdJ
CZbmBCy2noFYnC9g3BBF3OlQb4Sd+XUASUwPaxjtW5UrORgyDd/QJLQa3KPNBMg1rLT/uFoxKY8+
zL4/clAGlV9S/hFqcOllWgczKhDreLl+0gUSCwBZn+WB1wxLgTofO7/yMJv6cDPbd4EPicd55Ts9
7DEQcoO5xY1UDuabjXr37x/3DOn93QpMBrfbz/bhBVcGMpE5+t0dVbf/xG8JVqiT2hK0Kw/AlIN5
qjXv5RWBckzYoaYXkJctfmN2FMmV6PfFB8z0KMj7KuxhK33I2CqPFXTKdRj66km3dUu561aKSQiI
L07Nw90JUQsfAZbLdyDgw3qe9wyWBLpkqVDBptEcf9xItjTOiaAwmMns7d6KDhmx7t9sS1pmZN8J
/sgMqvpXjKo7wKeTOo2gaTNRIdrn+YC+mlGMcPhSK7Jb/QxY30+Et3saQF57HgOJo6SAjWEZ0T4Q
PDycV11pkz6TS4TGncQIinr3JAteIzTDS4ki9wu/LukkyScrgzQYeCJAok5O+MwNTlfOxXV/3XA7
yupZHcKO7YcSxAbJRpzcjowwbbALfncc9/0OwcSqEwvMG59ceXchNUptFOKRTfXkjVbZ919FVfsG
OlljqpJ9ASHNOx2FT3ZIUgkmO4TOKZaqqWTtmcAXpgxxUQ1X/MQI8y6sb4du8nX+Af+hCy/aWs9O
kLQfj8oKCo/ve6BBkZXpYOT4deixgmir0SMsgm3QdwOBkt3ldLReolFPiAJuEzEa3s89qKnDiizO
EzTq68LGs5yE0xN05vKNYLOeFMNu0YRF+A84u7nSJYia0/lxhfwAcoDo/ziqmDHAA1Wf41dfb5bC
gt5gjHMVs6+T7JGEhDlGhyzkRnB9nuR+XImRi1iOkVVAQKtxd0R6Hl5kxzQT33kPQXfgJP7kLhlS
JsS2fE1HKiuA5/TxCqxg3aPrpfBDunNXCFiR+oiSZv7cnVeyoOFf2oKkvDEzkEFD7NsrPWpPRDKZ
/ICsMzhfMO6PSiS80clHrIZd53b2zRud9E/AmhtAdbaYcxGoOlGwOJqlqrVF67Li6NrKV0Ph9c7P
s962gsFRR9CEkaz9jtBwMyIumcdG9ve+c7vTvXI3knw2OnIaBAsLwdNwR5L04BqKrShwPB35ukeo
r8dvjTR4e4s+HIJj15hEte4Xnh2tjztuhdCs0pQCzd41UYyFqEGxNJT/3H5ZmgSkSEG9g9ACrNA+
qmv9m5m9crgeVlN9Ph9rMkyCv+t6S3Bi9sh5peV+oHYU5E6LQwUl0PU837jF/afpslJrnC20VOfk
zBOKEEmo5uPw/DdCQGlmHHwQ2Uxgdg6T9Ym0klVr7ohe+2ovaSJKzHeX+L0rmIsKzQcAY+m4QRET
QdZNI3sRt3OQcxbJL2hxrHg+R/i4qMv5Swu+pPSL6xLljZrgiTH1Uh8ez6toMKymHdk5PoQv/YN8
kwEoRZKRZWJJhDM5VbEQHT+Hd83mBOYDr6D0DKCpKZ9E6e0RtHCileeS1fjt3pVa2UeUxw3e0hzr
QGuTl4GBxodhi8ktCAry8qghkVSS6Tg7eFvgGmqP0HdJqUvbXJFZsTflCPenzhBosCITUy/QiEMm
YwdPH7j8zPsDM6ImhqjeseeVipaz/bUtSZszKmSLmAO1sGPAn1ms7B4HYkzj6bzkPKspC3n91CGn
ybWo4eN7GZSYmMJkMZzn3tl5L4WGD7h7z5aMGiRWWGERnM9Pri1gJbKUnjXV1Eh0xlQA61vCCmHM
ASNdj1O3o7W+NQRhM9xm2NQADSEgrEzuRgPoFYkf9S8nsUzzKIhIjkApR6xJ+idq56mL4HqnVSPx
um9zEqfVHXC/aTFpLvKjLEF51PCctZaag0gaZ00tNBFMsp5Qf6rSiesLKoYbQlRad2rivuiJllm9
UyByhyUgxlplFYcP9y3bG5FU6ZwIGKG7oxsnAJx3MVqQq3kuaCNkkW4UCSUtmNT66V57wVQYhVrb
9AnmLtdNXqY8UASSF1R5woD2StrsMO4B6tTGfNHKXdsRqbMSLAPhzo6f8j0n0MYscyWpI/i0rohh
UDqVDOCk1EiTCY3CSpkLNT9qEhZht4e8zJrarWsnMMaIa6wt+RsyfiEJK+C9LunDOeSeCC+nElPX
0QoEF/n+TooFjMAjAafgrwjM5I7inIZfNhtu2T77ZhViBKeh0lD249PX3ebXq4oVBd+n3blIAvq1
If/z4FoV/jRGFrLroFIUUrmUgns4NY06/vykOQ9vipoV+siKFPzxuOcA1GTSdan//KSit5pjoGEn
5y2KFUfgtXEs3Ir9iwCiUVXJyf7ngiODtGwcfKexRal/lvwF7APYWiwomv+vOAV/A2pyEIwVLLqz
7jExrn5Ku6d1uqKIEeVuoyFOakvyAsBguYn3GIer1R7IFSrYfbW/GpjLrVjXSQqX5ZNhBFzm7AtO
WIHsApopr/TAm1BP77LHRRSNzBfw1SycANlLPEqBkJnHISXBFVuP+Uhx0XCCd1q8bw2Q5Tpmkb4+
p7T3LYIPis63bkkYW8AkoEHOamyrgDp7XxiiYX3vv5kngYpKVRdUHP8npUB2K7XH7LAXDTMahQcO
LE08NqOha8is761rC9kYX3YIwGPEBqNPOmk5we2hSGsYR4El7ysAb/ziR5XhrVRdfAURqKVnj/CC
EQlwtW01CHFI0T+PnLkJo7z7M8SXHcjrk2Od8Qh7E0AMHXJbU/CB4A1L8scMM5dFVtcbtD80ZY4E
Xlg/Me3bHVoQn/qO+joxIs9zu++MXwZSl4WeG/lT71JqHR70wqP0aQy2Z+l4FeyLdx96D+kCj0bT
VO7kKTKJjHwkoZmgJT7CE28PpbASBpFqbMHlmbMuBSBjsxCP6bd7U18qjnNo31ILZNHhPZR7Y8YF
J7Tly3qLP6zrF+k3w3xw6pa8oKKEoS/0Ed3F7ArIWOCG+danTN48jpKvQIgaa3WP+Ovikr8f8jHg
kAQvy1StIKKAn43QoAzVCEuLU/oHWSnqHEU1QtXSAOtL3zaonavSjNJLqmxZYRorogwrO9NUrStZ
Vt68gjA2e1w+sXqR8jshGBFUVdckOjdcLvHI0hY0shPh6EHC/MzuQmfGaoeSsTq3jrnl4HcxWFl+
8gMMLQYhgtywWMwDUaxZ5Q+CwEqaKpv+7X+FGKEUT8mAzzHQxoqPcbgJMyFwXtV4vzk3wnawKQzm
UkTydHn9NxwGQ1PIXdCnIMxb8srUyOVM6YhloDicXJxE0TzOLuSEXYIrgpxpbrFofTCQ7D81AgBb
BT1egKUwjQ6byZlv+6xDMQwiNj8yfK+KPsr8Su0CryUxnHQNDs8BUepNMnBRZ2TQFRxNStFeNtFR
YJrHwtK5PPoEB8wiElC80+BO+xQm+pyj3vgh23aOVaRIvUUIff/m1TGOCUMOCNiGByo4fjbC1c/F
Bv1TquCPeB7a8uQ+DsVyPPWaTJ5nbeK27Kw1Zr13JTZN3eBNpneP92PwU9QHbYPqdfRhwd7dJVbD
I+SqZKzTYu96KeF/jpyFIwciIcAvkNtTheBl5YlYhjDAYWewwnYOGuvY9VJt6P5U4bs16YmwWclE
Cck5bNGlcV2//p5BZUVEDvZEdB2+cZDf6npDZzh+LM0bi/+PnCcYR6naY8jxNPckj2107CasjuRu
Ge2x60AY6D/OV5RGIIbR+MgxDp1nr0CRdiFLEaDk368f4xBNgAJG3fGkzJrfNlNns9vYU+wokHS0
14GJBeQcT/hgR/EF5GsYccs8/nPmr+ZygbUPg1oiBTvHr2itkCxKKXYuEdoeGsTnc6ZHg4xsaTaN
Cg+XvXxwqpfNE4DXwXFiAuHtIeZpFF8ZE1pFzCup6uAmaSDlgRyc/J+9FK4nwwOSP/+euk0zDMOP
ll3rWnNqWwox812UIoMH7KaT7eTvhPSH0ESRIdZZRxmdvf4tgGt+IzaS9Ctw86OQJFo6XV7BEyDJ
zuRshpBQT5sb0BslZQCJTByTaPXK2Ckzt2QzZlt7fMTsuMPV3lxXlosv79hpmNl27ztERq7jjszB
VY4TjeoaD27WLmATY9qdzLY890fofCiasQKaNFrN0Bq1rmX3MDg2URLHXjr+hWrEIeR07sDOiab8
ShlCuJnLzTD+TMHzrhiE1JlYCQBwt4ZS2vi+qRmLYhaq/ZPZ9CpkJmMcDySl83rigA47x/8S/0Dy
3u6srGI7I9kjLENVgOO59/pVwtS6MkS+mwKyULwKJlMnCqIlEHvvdZSKnqhKZNNHPy62lV1PsoQ6
LXDEXuWCqiaLbVrG6zELw6yWpVKwOYhpj3CggU0HbUBqPstciVtCeluETVT+tfu6Ju/mP73EM3Re
j9H4f4V4/EEojbNwH33LaCNFzfxva9u3RTt1i3R/zx7kt3wldt0egGLGNxtguFCaxWXuqsAvq0uM
JJyGb8EgtN4VF7tTz584FXwJXFPuZ3dllqdm7rL7zSjJf4QGdaeoZqIB1Kpeqxxt2PBoUbAFOSwj
hcKP5oIWTsUElBThR8eLI8W5qqDNJg2u/3H8n4sJ8BtyZKl0B4UiMu8eyu0m9yqo5Z8FEbSMS7nX
CIsp6o6SDitybHEaKMoTSVby04+RLQVousFaaPwvLTgTSYatg6fWga3fKBSBcPAvjbaImGthONGf
cSk+nKkXxcmXsB4hrANykShhlM6//7Ebhz8h08uNEHDo2/dYuFye+l6B2gkQPMNw08KA5lRdLLVc
FUN2cKNPviivcII2leOTU1Xi8p+dDALZ1T6iA8EU5QGAv+AUb1fNga4dyEO6C96fUNknAUPBuzm4
oHD68/VgJPXYn8xbezwLdYvXSX51uMYc+NxKlrKYpCzk+dXQdzJTVozShunsnjTpXs0lO8hIUZpa
+O8A/Vf89VExCRx4+B7R4MpxV3YcAX9ebSGwTwOhNcAAFkA1A7PjBwMOG1cFtSUA3AjP/gjdXZyw
Uot1LWIlcmqdSHtE9WW0ZfwCnKACv1+9FnBjaeLSS0ubAcA4WigQJJGzp+uVAJ9W1CdqgJ9dm6Tw
rYmJjcoWq6OXUNKXRhwxajLOkv0D/9Z5o/JndDYHl3/l/8gLrLSpHLN+JNIyDV5awrUECaJpqo3T
VlVk1F2lvGuBK5wE9wIwa3w59jZYSXpyIrZJz8x1J4sAcNptbjkMfTo7j4FXJguEhhLXoXhPSatu
Ie3LGsh1356yMglmO+F9K4tm1nJGwhmy+Sn/HWZPWNMT05KuZ4OGnWMnrsu+4qVV30R7f+pHDHvx
Q8vuDZf4jzrY37b2P1W6Ouydp3UuFlQMcC+Y5lcMwIqDWL3iwKA57HRxFTo8FpLZwQECRWu3+Fzf
+Bi+SOzMFYgUzAl3mqCCej6IpMHl1zIsZnHqH5X6WP70HtGOHBmZc48HdeA+3xxcCK4PTxmxIb07
N8Tld0tlmmdXF+J84Otm3Iyj3BD4iSiWp6O6zbwzH2vi0IPCAu/3jIqAyojIQbMQAP8Tt3QUOdgn
RkLicnsw7+Ll0CCulb7nshk1S4SW4blNQzsIoAFl63IfhACp7H+gRjT47yVcNOXt9moFUab83YPN
EiwtUzmwkBHg2u6cjlCcKsPGLwWbarCupiabkQy6wO0iEhNCH494JwAiDklvVFeo+iHRWc7xy87p
9zXwSYTvdUKF+cg3mTCm/Cm60lA4GpdAwz70YIfUslrkN2YtQbbpvHlUXM0oeFU5oc2dGjp2eqZf
jwMe8xJQxoHvQv1zTYVsSWGjFtpdikFugVEeJNU0vlz9f5L0pLELaicA7dO6aQ0OMRyGbKlPUEmI
1Da8EBLVxAN0SJRj5sBv4gLei1VkAG7b7YzLCyqRpk3iUhEL1/Cq00mw5f+5VYl8PhA8kH9z/iMx
KycWduFPfNZYY4cBX3SQcJuiv2p6OEWTdsopSX3D2zz6CkxOME7ai2z/eLed1fjKfgOI2P76fe2Y
3mrZ0/h92SuJDdEk6YVv+WW/N2LlYx2HB9tski/ayJmp3OiLqAwk52WDBVQgnI1EtVpsLN5RYiAZ
te4nHeGCAO+OqmkkzZ/P0Gmervl9RsxdGtZP2Ue4k2OJoO9DdSKR6VKmLudikCFDBmOJ+q2VL/lg
hY33mE89XiMGKY4GWe8FJBm40HklN6uQz2WAC6vS+ILl5nbIvR+8g7kZ0MrL73+XqQa4CItyWoqd
c1N0jpp0EHmpAri3vha+yklJT0d7aYuvGyPWn3FiVY2vBArejtXyyGcL3ZwV/BFjhRRmtUeNtOIT
bO1c2/wI18EIv0h4SbXe0zqWqPRmGF8P2BTJSCQja4HxLi2984fM5q6m30PNc1+3PhfyjPJ9AR6S
yPuZIziy9WKJf26JVNe6ZGas/WNeK+q0nBu/BeEWF1W+g0a1Cbx1ondU9JhvxfBffkG4jmBdfujg
Aeo1/umGr7/PGa7oFIzBoCHadDrA+80G6HFrXF3e+ZLEvl+Sh7LPoHVqNV37G1ptGtqcehLvZP+B
P3k4lmSsoMWXFz5q5VW30UM3uZRg83JZ1BUf3uozSb2IwJPsuNw1neNDbF08rIigJNP9Msj75+Ke
C2pC0tgyKFPrL7ORjSsmLSYOKaoXUp5hGMCRmiBPS32KWpOCfRpZOic1OSmaHzwKUWtaLbrEhJJi
mqH8y20zbhqPc4qF/w/pqhkMgE/9T1AYvexnJjLKAImxvu/IxoTfrRRtB+uF0aXFHaRIQHn3h1rK
YkUhmxRw7eAunaUVGW1Vt+aUXAKvE+PTPae+MKc096aQsyh9bGCiCJhePzYGq61OlnEaNYBm83TI
wjYE/9uWRQVmOio+9g/QoYBcz4Ul9VTs0/NtHso7nCUna+wh20VIVNZWfzAPv6BQT+LvsOQITzM8
sjf2tvVJrrMCbFzGU1PzMrIRdX76lyLGBuxYkPgfb72Y0iPVnc+JLRZYi6uc4DYOLiVOp1htCa5j
nypb9x8b8toztZGQy9foK5ThQ41rxgXl/zwcs+nsWTDja4bE0uqj3IF+5gOwu0YX5P+GWF6R7RUa
JVMeOHCJee+2nr1v+OLl/OD0DfyHZ09rZsDHrGyCKAEoPOoncEYO4iIxRuzm/QgRTHMcdx38nhwo
qPBOa5XfOdW+ZRrn7cHcyna5NSOfeglvXJKY8VlZlcegjThgC/6M7TrQkaYk5GYTmw5pusRjKAF4
094kn3khYSw1BOD0ygNTgvfpc0MseECJ7zirUN2kJroFJt/kiSkjxKFxMhYNT2FimIGHBmbTSyKk
USdKo3hEIJYTcp/dx5bgAAwfr6ux0f1GBrXnpOKHjZvrd1l0StFKA/Tn+6eyc8O6kamHAzGOkHU5
jfkMeZFngqcKw4EWo82r1aB/a2myqH463Jg3UKfTUHwEsrG9a5tYxVqeldVBkSoXslKobnYm5AqZ
mZ7a0Uox31OlIHhlmKcchd+Klb5Tw6Zrlw/8rF29thzE9s4gCmhkslhUnTBIuB6ymDoGz1q0NBqZ
l3UGEYR7HiGdZeos93ismYtCimpzKTUZ27kRtE0tI8d4OxgTEPp4VEF0yaEVXPf7bur/SYDvSH9k
Fgh9qyMDuEXmA/1DSPNl1e3Yf4r5InGOvQ8Oe8If+wRAznPDsdDxcdtaKY1Sq+FnQnDgnYCsXVSb
MLCq4gGs/YI5uiET+GzaumKTDv0J7AmPs6DAT26z+HHMMmCcCFZt/zCuOQsstegRxWMooQmuCLpF
rnNhiRsOTTAZslOWEMzESw4BgrU0Mx1QJbx2DN0eJm/s3Nj7UHCEg9GuYEMUGDdu8JkBLqILXbVd
ScIj+KlYVujGQr9XN1mVuTMeAlxg5ZPcJG1TenrlfuKBq9P1aeUrsPvWyUrBx4Sx4Gehjfc9Sm+o
aYBJukI2gL2XspOqSZ0l42zySmkVVH8UIucjF+hq5x7uOnYPh+azuw387D58+Qa1Hkk3fQnzvjsn
e3nb32cbKZBEFgfN6VdCPL0d5hwXFb64sNC6didSxOYyBXWDIqAdsI7aYD37hvUhLdlK9lQFU3Xe
muA8E3vX+aXu960wg9V0zni+3nkMVSdFHrU2lF78a6upVMWfSs4xuoTAW72Ex9QeIh+H/MUnUzgR
XC/R2f0GnWN+WVMXDipIbWCVYgd2xeo2vyginpnE4FEk8b8GDcrE4pTJFyJARIFkUlpUM88836cm
CrrEuu1zMC9B1PUDeALgy5MLe9fK7nmaqn0MS3tfDvKrjXNFji+n+cP5SLW0EqPkZCdc/PnYNfEt
Q9fdv4ykSWizu2LOYaSLScy7d2iuNuFiseBhSGI9elzUnqXUBAlvmFaOgsv794c3tHv5tol6bF9U
q2NrjB85glaHI9aAeDrzcQB2a0ig7dNaYEQCNy8o52T7Ld2Z6aX6RgM6I6XOPfc2fq79+EpPSmeZ
N8YaKDicS52dO1s8oncpi57ZxDF36bCW+jf/loPcTPcLd0IcxwP/6WQ04JPiH1saj0FIDL7Un4rR
zhm+hYHzmlMjl385fAIfJ6mIwdysCkqJ/8iZMfBbQ8dgrIQogTxKTUp1HwXCBp5MVUBCNidGgZwO
lhVCeVz98dsgzadUnshDQ5NrA93zUUyfTBZbgBDPT02icl8qN/mNQht78yVWBubW7B1aoX+0k/fe
sDOs1L9LenwXPI2HsxrDuUf9H3ADl0h5I13Gx/YZK6+3t0yU7CqEPwnQIL4dweMiMerBWBTczE30
wy1XycNB0dMyC4+1w94n0OcdWlrQN9wN58FbWzsEk/LCVvOt8yeTnmcXTbTTo2ld33jIKItvawWb
sLvfI052tfOFEt+cepvtoOCJAeaSzaGbb0daE7zvvLQasSnGx2i7HtbfzNJk5PIfbnrmok2wa65c
Z6yVF4x51psZ8VXv2WHAY9yiv4AkHhVPWiFVDR0zwmGs3/Ljwij9h13jpxQd/nQdhjq1mIF2uicz
OBqkgrqMbgoUxlvIIz4TSpToaa0pgwuOMYZ9uVeO4RJ9dveI33atl9VpUo9vGb+beZULYot+52JR
33+oUU/UzoVDtMwSm+Ii8gqGRM8EI72zEj8cj3UINsdSmO08YhM6hK2xZ72KPUI0QXDEweKzWR0y
JZLbV9wWFs3358wVTJEmqWtm7iNjPjTiFjy1dX5TG+CLaDVl4fLTq12t//tm7OQ9t35q12IIuVJ4
YDIEKquvVRSO1Ri3dErmcQgF8bQ4sfVCOHXl5V6QOzDlbwaTgZY78n3aN7Hx9vmLwQGCECh/2t3J
X+kBtEX/qMIpb59l6++n90ptVb5yKPVh0ooofMVpxjcYuffKQExyMQHpZxFaMHb1NJFyRftlDbRJ
a9OW/RbLaOal6w4t+Fxp+aGfrL1kuAKY2bNM+JupcVRsxfNRzMZFPhzNhFZaM3smokl0PHfMpUcg
/q3AtvCxe0F0Hxb4lczXVsQCiHxG3IszA2jQ5C/+zlNEYD7Dw6bBSqaEMlS+2y3V6El4JG+ov9X0
NY7BsfN9v/DliKu4uArkjE8aHlA6UzGYCc7gn58YvpisPrXsotZ+K/R9lvcve24SaS+0QXbSnrjI
9SkXKhRShD0mzODL/ao//FikPz9/eMH5KdwZIjR+5agtTgD1t9xHv2KQnKSD+5gRLUNMwIIgK0wF
lQ68Q+oT1HZzZZIroJfS7kdqY/dfn15iSBT6vTN3akLJD54ucrrs5pBXggulKizEEpDL86ICWQVe
vUDZ4JBlek1ELElte2dXVv5ymhhDAqvSnL1lzEp6GlYWI6QFX4MYNvH7NVJqdJtP2oWZYwqqCspy
3Uzcy21gCdZ6GGcXfX1rTHqf19liNZnsBRbmEP95bShcVBKKENVebNa8CzDgcROQmWiln0gdh2kX
wYAS73VLCR2YX4ptmXBoAvAwaEHvXTuH0eMzBQgZT4ltclXkcLoGrDJP0M7Gwr28GVFp3hbs397y
+w/39MtwTyLI5GxN56cY8GBy9VYGuslwJGR0wx2BVsJPI9PYDouNnFfPcrRtUsLCAkKpRUtmBxjm
I5ftDuu0yVrvyKCoOZOr9AB7MwN/MI8admSxokSuta89KKxGNCDuC3mX3bNrseDUD2hKAfRaIvbh
dAkPDOu7w/Rs9kt1qw77mpMS5dP4D2GQ00CUyLu7i26LmnsqVY1XqyIvSo32Po+Z8RIZJKMQ/r4A
GVNNUtJbC1GcZ7e7MUm/6cYXSswCfniuir4+RV5lgc2GAZmB3Ci+F1owo/xjqk7oQ+4Fl7YCKL6c
jWprI74JE0VdnDc+LCreCDQzLG49KwyYiT3DgplU0OSXJdcWSVOeVGM5pVrKkGWGOcGbGo5FaBKH
ebACOq/T88Fl2N7rlzensnHNsd4CuwugCA+OvY3Vryu1S1CNa2roiIbtakDagCf72W16sNhIvv/E
CO8aA0ANIkMs8Wk8vD/2ozYQXhaFePIHl2ukcFAPS7AvpMCB1jF4/rT9ydiCc1rT4GqN2L6gxjnY
TQLvOmqUJeHmOZ+GAvkjbMl8KlrSEP1NrsH9RQYXd+Cu1jAmThWD9ExYAVhGVNwHI73DdLoY45oG
m+nfQZXoPiaPuQIru6FnLud+3YLycAw2lskRkp1cVNb5cg0a5ZwYneEBDk/ZGJhPGWhDZN28+iMT
DJTw5EZq+WDzU0eT0isAl6zKbNCJNNVKVQ8dUSYnQjSB+7XSwv5FCylOsl1tGqkYW0o4MzoI9rOt
Qkb1zNIxtjV4hjcko/Bipg+BeZ6LS9NsLr6Otr7w4apFUFQvRz3p6Eh9bau3cpgiuCKK455v/3qw
pEDGXMFXTxGUg3KjuuAwvrodxgLgNypYjKAx2YjEnmRky1sXA8mJEKr90HK5Vgz37MyHyB6X83Mk
jd4LHbR7ki9PsNu1lSzS43cpuiSl5AJHGlyqcXyDjQQUgQvTRLx//4b78msdMCmmBzyOaFrhPoBq
cJC6MibpfXMZqDRx+IsfvO1Z5xf8EE3Z2VbGaXhr9S1Z1lv4WYIby83u5+d00UiIywhb30mCLQSt
SZLLMkjbrc6gnieFSFnyUCme3dmScwqeBr0W6t7fqQhfjWvE2VVpxnxJ5gJs6hTznpq/F+L+/NRL
valHSmcTNLJak8e6mdvS2vocfLbA2jBrmu9i4LY7D9lJk9fOoADIpm5H9+75wYfu1Zp8Sh4MygZA
IVSvZmnnEDk9LP+gZpRR/5rXJHDjm3K9r/6mGwdASUbuoV5bRIWli3puwxfsl/ANnBt7ndhy5DV0
lhxTloZKSobA+jdFojFM4TQt+Ixuamdeu/IOj6Q9t87l8IvyBf38BobHE/cEZPtH2Ja942sBqPtM
3TfzmMB0BnlWR/q2m9zXcyW/9X87e9hpQyzrQQEkk7DunLugXKaOUjcLPuZcuXZs46aA1BtL6fjH
wQWSM75NNr3NKYi00Fz1TQIIghqpfDN77/gr8ytx4I6RkOCP5Pg5SSyJ3Yb736lCZQUDStaAHRHc
f8/tmnI355w4wJzyx9Lw+5ueoD0P/S+n4SHRdBJGiMXnrTZC2p4lc7hF9apqqiJldwxF/3e8FBWB
CBoLHavoH+n3M8mLKYZv7qWsjttutpdKwBpUIdFW9RPjaBBd1TuxgAxQVJJG2bSyVSJmEyPB1kWj
F59NpNY643AoJE34RFgZjUIUa8LBZQxiHJUmo2195Cs3p1vCr0Ma7TE6gyw4aElRUZ95lJJPdVKN
vV727xl44LqjKX204cXjMAIdLii+lg5QAnBFWXOQM8OjVPjukhScI9xQagm8R3npVXRlbGAII7Qk
Uc9sC04AlmHgkq0fbh2AYbj0irNWFDiFnlVEDbiuVACFHBHIi8p0FT7pKDhB6rXWZxotKQ9LS113
EkEJWohshDv6aF9ouaybNgvAQvB893kg2BYZFLE+u5+Zm6w4rUsVfMjn040sT4x1R0L316N1LQkP
CSSl76SGvUlTRB0h5iXhogtOsegwu1L0TXFKiSfyXI7qS0diEXMPHO3VIFg8EaLZwdMv54q6YOGl
HBLoVa9g8WdT2w63f7hr5RQaxFP+FJTjcZiiqUjdJFopg88e5K+QdoudxaS3lr1Cs+MrUby5HsAk
Lt+gvCAJ2Ke9wU8ou79wAShuwrGvvu38ccnrmaqTtLXD0ITUwvpinOUh386IjXs0XBoxmqHSQq04
bTaT0X0jm1bLrdzRW2Caxhh1hbkfY4AVNaXqBqYpKYTtjHcpRJMImSXfVj6Sdy05k6FzAPQt2DKb
ap1npX9ealIKDUfmMeiS30f/y+DvgnFmv8/5ctCALGT+/Cbs7S1FaC4QElCalnGl+2wxBHhimu3q
3TZDdGHCGR3iZOzXHSLRZu9jGfdJUIhsrrUAkBqIOPz1VJYZzeNVi9zMxH5xLdF0Xq4s2EphgDI+
LSogQWOMYh1Jzii9AIfQvyfIlTw8RDznOSEQbBuM2tC4NxmUBBVBf7fqyG1oQ+NtPxXuNMaIIHGq
mzq7XxxBnBJAZmLaZQKh5gMsFV60N6hWh82+eXHtofiUcsyYiEicyu24jBNGNc3D2avCoNonx3HC
6Hyayf73rPreCD3wKiTSzfTKI05GWPSXV4A3ayGIYNsQPtZlINxe+RcBbzr4TJbjKcCWALTQxcIi
wa/bzuwCODW3jo2yjjj22sZzxU8I3EeFhlViTfjUxzCcwB3MOuUWaPuEi+9sFBjFVgFqdLYUMWIt
N2mq4i8LbaUivbhXqEMtSBPhYNPpNnGJwvNTmLazo0OIGjeM5tqpI9DwEGTJjCeasTxWVpGcSIUR
bVAF6QpBi3FjnYOoslWq7uWsbq1gyqkP2X8npLAtUmynB6iXj6xGAVZsm3OB3wVS3QEs2WDysX7F
q4mML4Ahe16PUQ7ZSyAx3WBirBYpASkmJPgX6/svdGFhSSiNWVmjBmMlVBBQ0T8/in+3ZZY+75bB
JC6wmCcmOHAIB8o072fkzcYR4KWRXLlF3YpZxrLe/UFJnp86PSU+tKFMXSTbtyY2Mp/cos2JyeJ5
R6eHOdOtck1WIrAxKirCYqq9WZykf/ZFD6wAXrdmTrc1hQxJWMNZwy9Wc4q1eaYCve84WucA1rfF
xSoM10cmtGN0/ObmZicrIO05SjXwj9Zl4Z8tE0/pDmkandzRKjUkQ+RRanfHtY7bcS0bM1d+cT4r
5Usx2SHbV0onlew64PlwQxUdfNnrfeqBWhiJWKj8ygdEIR0CQO3zFGD5ZmM3muMvI+dDMJJBejz1
2LW1O6QjvkdAPN3vwZHgQE23QUyAUxlTcYWeiqNHVhA4CgmaYRR4yeSPbUeO/3DUj0ZlDiVGbCeR
R4NviE/0Lo110vBkwv7DT0jfuiaa3BVXi+rk76jAvixXln4PciR72z/V31SRJE36IaQ8JQhdlq/i
5SdWlUgpAJYoMWQ/AQo5saM54CIklnrYWnxZjuAslAWndWd3ofGoA1Z7QzMbgvo5a3egB0uKOj6Q
NokO4POeYQXyHRwW8AY91hnvAfpPGkGXIuAKtdzccDZvPlCDNV2caKU+vEzkG/VjdSIffJzgyjJK
HBFBe/TAgWNDe2g5S2z+HFfd8zb76OcFvjLbIMx00XL3ZazH4lu32ZvFGVLE7mN0u8wvH51tkdLH
qNroiJ58nDAphterm0tv/bR2FxcOjYQRJHalNmMHzrUEfbs2c0rSlFUyjysQt5E/pjW/G1WglJdR
Jq57Q8/VE0UMaU+JKa0GDC7/1I6RsHOyjC9/ChXd7L5Gc0uRrm1XQgJYOMgI0+BYpB1mQh4yxsnD
X+fvhcRwrpzfR5a95/sNL55jEfqXknI+Y/4V9D5OqZI7GrgrgPHba69XFD+cb8XGeV5PatiJ4vlX
l64mC6UTMwtvlgX+oKETFE5RsftLkpqythVb+1CX30wWP+6OV1fII5eJfFN2CT3BtnHru77uKHS5
pYzXuFQ6xocyERDnp7CpQ4IDcsf1gmjEY59zL+u3kepw4bLDG3pON7n3RMAaooM2+rBPt8QLPf+h
ZfT0Uz7+SXI+dnHwVKOFkx+AxOsJL7DxpwZjF7cfIHq/AFX4X5T094hB8rEDPAGG3ErWqeQhQ81X
xKkLrcxO6UityXkl0tjcKqt4C5yoWUjAJp0Q12QxHu6/OkukHIMDYAhXdI3galxj9khEMfxipVmn
8PRz+WQnmnyDrW3OEbNWA5+rr84UNTIOyunDQ7qszRcdJi/NilKsy4s11O+2787OHovvdsN+fAMF
kV0zvxm6/clV5xMY9B9lVJ4R9E6YR3RMF6QJsISNVdMjJrB/kpQ7YETPshzLgQl4l7yR+/hbSwkr
JLqGdYxFGW8zcDj1a60yLJ8F0YY/iA8HzA+DVOXitGpWhmEtc9ieiJAPyr6J9GD0qDu8QCHT3ePv
wQw2yO2FYhzN7zmrLrjA8LBGH9LmBS3qsedpdiSbQU1jK3PzwomqKh0kE6x6OAloYBHgfEfsxaqO
4bofnC+CbNpB0AyHODoYvp+oLUG4NN8oCfRXDDl0Fm7uorRW9GI6cHXs7z5hssHi44OS6Tsf7eS8
OG4A7Nv6d53T/1COvr7CFbCr/+ZlJ92Or7L3kdWpYCZmvuaB/MLqcEzln3dRUM9P7nfZehx0OXvY
x7ZG2JPBvW5MFefLhUmoWsZ5IR0ki8SeqefTpUbWyE7qMKvHrixGVQ/nkfqWRQ28bgUF71mmGqrf
MqafxF0sDQV/HHtDhTV8bfEe8lXIotUIMABCpyx6kKHlzBTJzzaTc2u4N1RulJWlbX0kgYYeFRJe
oeYx73brFc1KsUnq+KRnm9RWYaqkNP9G9fsFphXNAc3aTjMPVhfjMTTKAjlpu6rzee1qQhHbbrl8
8MMnv3xTh9WW4Jre8t4y2Rs9h2wNusmikH3+BRvoe+G1xlokO3GDJzE8RDwRok/SwX/gZ/iC5VXQ
ZIsZ9ag+JXtRz7w6KTmKurZG4T3IPWD0JNT+D7JsGxoLabLLucIoBSbbqdvzIg66SgLUWom7drbO
K6Q6fI3epa0fkTwjVNTIQ1QvEUo6ePFuyw/XvhwTE/b/VRWqNUJ+3dp1ABK1IoAullbgg95eqXPy
O1OGSwD05kr6JfG4sHI+MR3C1JtaewDTZiiAOLI0L4wXdc0poCeBm1Ip46zy225PO4LWfuMtjvYF
LI2+bFQ7gHCtqRKJq/6t/fuG4m1Nd0uncc8fVvRwg63dkxdGS8Hq5ek4vTXj7zQY/53F8DOuokQu
y7jHcFCqIUZVvbkfSxEjOAtz1E2coYXjEcYABtST2Abwxe+EC8KwQrYpJDahvoJAtsAvyht3MZdP
DIDmdP20xvwNlO1kbB2leb1n/IwbGbdZxTbC+UX1J29j61lYIm/TVLNm9ujDIKjQGxFTdkgB1Lie
OXm96H0sFkSfdFoFTsYAukVN9hArak6OdLDOdBo9S3xln9BpYzkVNKOggfDirwnysHRfj/W3Zuix
GW9woo1TIT6pLwP1kPkaJGrsCcrHBqQZxYAA61Rlq1EiWwTWzct8/1zct2z7lJ8tHvIDZKOq7iEI
JRFynWvCaP9qQaNuIDyyPrlPvkA5PfQp+CvaEcQ1uOUl0tVXPv8OyeABV+4TJ03H3q8fwpEFdAxJ
ZngO0/sJpdnZcRNM0mpBL+6wpTOaD+U9XSegv8z8qRzb92VM12GDD6k38KjdLOLqsQzjRBpH2JGy
0ymlcbVFlDtvFxMIGHYP1zHOxU4JNOEbWfC2F8Nr8jlpA5gDwlN87Clmp1AOsFk3J1f8bcmEGQja
pwOPCY/Omv02qhchMpVIs9DwL1VyL9H7LQf+PMRUZ4MycBuuncXCJJBKgRbvYKs4UHaBgMi78O9H
vv1HzgfYKCIIRrMerRksSln3ZRlJEjvdmycg5ayVLSTqHgeGVWyTD/5GUb5Hf2A5ikpFbbsaZ1d/
J0Ll8NZBleiiXBoA0oiBmQa4saBUhwJp9TaZHTwC3eHasY+aqt8cXgGa4g49Seq28U/0J1UnPfQW
Pdk06VN4XZg6+dasOgVqs3M3FHbqWE/caC4rWh53WLlMa1tO6fQPtCjwn6uck1FHpYzoXt5Bt8ch
ciU02hvOAwfNytXkYbQIanFSd73Voi0Tu3qhFAT3z/KrhpRoK7WsRO06VTkd5pMe4q5iOtGiUWhe
C2LoVzkAFhSOMLLQMzHohfqpeKm46bdUS05ZAxAw0dx5/ddOVTnnlYaoYefAdruOu3hkCfkuYAG6
zqo0rsn1Ku/8MPDEMUtgDRD7k9XHwDEfpKlA8JvK1K00zcBXGK8I8qLMlHWgXus7NICen0g+Rqk7
nfhi77sCVcGwg537acC1txXIAN0suDgnyYKisCf1eoz4nMBWjTipTser+3rVmsfjYcZRCPh98Z12
mR7hRm04cPSnExjum2xC0KoYqzByGywxyFeTFSX5IGj8TAk9kK0p2aqXCXVpPen9TTcLVDNGcTYm
uRQd5xYqG6aswkQdr9K0wav1FJQ+80bgkblLvv0O63Fxbfx9sqFxLmsf35SdJMXS4KsdONoKSzse
5xN2otZ8JbwhzgZeZRs66y7wkQAB1LHIlpx53d9oRQO5Jbwnwuu8XHq7NMimvnVIMxyaEaUYEX6Q
lH8poSw9IeWAbwMcxyXmBiRotkCe03y3BHV7btu0mgRsiwsDQQjdI/kZPFJEN42A1LO7UCOjnHsz
bL8dtMtZk8vcPcsr7adtXeh8/WZZEoh679jVTu1OH3tCaHrPTuuj8ip6S28acGJRVZAgD2knCVYB
rDWXbIVLFqNdCFmJ8V7u6prTkY5+0CNaMBoeLZoLJypg3E3rTcMWWI1FSUQ+urd7YnQf/IERWJ6O
Cjo9PvBqOeBXZcfyGUHCV152oyE2aFsQDOsACI9r10uipKf95x7wK2pHZLGjYRWmL0WFMrDcc56a
ORyK40J6M/wUN0sxuq9CCrKuSUSM/usNyJehCoUyFAS96vIiwpsZ4iXf1pZdZs/4ahoC4/AohybN
UC3MhmdJqI8UnguhukGD4yLQkXqT/fb3OURx5JYD5o7GTrZdL9F4VdLD61yXtsFS3/jByM2VpJpR
8YNHLeS7pSLtnw0eoL32ULKjuMEXxewz7GX8Dkaw4+wNK94z18v6orV2d+F6HupTp8oc2xGiUUMy
2WKyJSV12yYkbdtQxhjS/w7W8yueHKm94R78w8rQA5ibWK0VIFGEeKXEY+o6CdNHnhQbxk4v0UUw
amP51VSgLHef7htzfVDzMlb3XDEoqA0JoWLhtETfZLGSvkbU40jteByw0DFktqc/wbzsaj7inbIp
GqvAp7qud7GhFR5v7+rJ1eEqRZJgG55CU5cagmDn8KOeM7XZn0jjJRP84Gpj9QL0Vis1hhbhXsjw
ckMFiHD9sDkWU+xe7xESJuVeqM35is6kBkQFzudkprp4wCXe6dsvglwLa92EQvSI73I9XXYdSBh5
F5labMUKHhjaLNU6V6BjE04ozxdiohBpggVTxOITlumU0mqKceNjYneYzeJ8+NSr6x+myHtrnl5X
b6LCWOEiG7pjG7WiIhLEwpET4ObIBp2YWlh2ftZdGphXDGB6TbrFApp8AqX3Wn/1n7265wsvFcuP
S3D+jTnTt2hMcBCIhE1F+/Co0vJttqwxWYGgEIv4B/mD0ahaSvd4Gij5e47a5yVSqVjwu6AKfb0n
yIIiTXFhNU9PG27SLilUyuK6/9fgdU7xrxJF03ljo1XV5z9UHkZUgZEths1xSw3zaFcb1Z5+kq97
KhoKGRBrDjT2Cmm6+92RPaOt2Xrgnq7DN+PthDXGWZ4GP8aPuAn25/hS02KQpSs35KwWh3H9YGji
oteV6ABNgjkY8XdmiaUu0O3tkljZOcuh4U0UPXzll26TnNgded+NstA4vB6bV16gbLJAAdlEMV0s
7NJV4MUO6uROKaRF3zD83S8/UnNlYOOAQRBSbW2xWgmn0vtjIUuRYoYarRjnB2/ZZ2GGoEg72l1U
P80MWKsfEJHgzeRQIC5rlyvisCtSHnonTW6EaobAvJ1nkgnLEq6dWES7zVhYW6kq3JoAfkKpOJOY
x3gPjSlcfoT6DUOXcOjafYGpPKt/lgVeHvQB9evsXQJN6XPTfPc7mEDobDTXt1kRlPA6xsPIhJLG
xIjnHe1qz2bGFBtcZ9Hc2gs73W49OAf04IqEyGs2q94gRpSPa02PHruNS1UMer1BWKPp/RMU8s+D
kwi9yn+JRj2rAHxG+dqm5mBzgFdYwhC6DoXEJ3lD/glcBB1hHJjnMrssLz94MgFCBhY6437tGElx
Yw0IUUjA7JtQlsCiwL+eXDr3m8YE0+ek1SR2/dYUsyt9Yzqug4O6HRWSsKPskvgNusxF88lRMiHc
9IooawDHPHzrHLZ3LfUSd1eoUNAscvBnE8RCjRP9VVb7LN9TLUPMM5IgirRe5F6UfWEmRWk8uYob
sXRcjnyPfVqG4RSg48E4kLjvG/rK+nNEYCSN4f61+diePLP17PYd80gOOxFTqGxR7BU6JrXlAdnc
ZpEqoBytqajl3i61eln1Qu9ZvzsHcKyUxIRVg26n2g8o+cPj6oKhVm9DI92Ij/vc5RscOaMvWH8V
Bi9eV1Vz8LdffAxLq6Ne44wfevoPuNokqY0DcroeZ8FYzru0TMolvefZPCoX9yA4i77ENsDMp1gN
7TPyR63p4Z//ydPCp6Sj4eRBicAJ081bFHZ6NuzCGjC9KypUkEVBcSIj1ms6VXRW+E8Dof/b491L
FIPxrUboq0fpKkbscZEWhMYsAnZFeVhdsYkpNpHzewciqQ2R3LCAZy1LBEXrdWyfdHu6XEUph0b/
Yg/8wXS93Xije55P1RxyQz8U/tmIJmDPR0ozvilwX0LLaySfogqmgFwHTtjze8DK3U0zukyg8kzl
oTQLU5OzIuR0Zcdyn6XZJaHYE46DOIBveTT8OduwcrxPyFykD0xGDtUu9Df6jOnWaN7m55uFMknE
sn69WR+w+0fjKiu4awPf/eiWLdPcIwyg7EecUBsaYLNWddMWd7PHOHRMnEmv1xGVaZCtyTUIMcst
tk3xGdPxGvbwbuG3zTvhaT3H5l6vfIxSdYYZDDv7jkTOu/pZLc7Ya/wCy3uJwJyrVh6tHLCsWnmY
59y4xO22ldRxDK9qZXdCGbziRxsUaC1ztZr/MQw/S01Mppp+N2RZ9zw1NvpmJ5/g4zpf9N1HE5GZ
+Z8H5LrGFpe0hc2lCiUxcoAqwoCASOlndMeKvh3EWAJnMDgDZ4R2oN7/S51l0vRtyJBtOb8gL2fu
5j679ZDNl+6nFT7GwwekrGP4//Vf4Nf0pyTYnOof6lt0KIiFcl9ggeUFw2yomJMH9SOrSiQT07yj
JpbyfNP1Ixd2KJ4S2FQENsX39ZHZzb5luf2jPXrKG2dySZBFacJqdLKNEQ24ALrudrqbsDUUjArd
zir/MG6OUScWpxdeAawCePI3c3L3JBQC2krX3xhhPD83d+JOxaffJn5+p71fBgx/sCzAhwMWMlMm
hX2vW/pk13upgJezpCzQZsMBZt1vaBmgUowU6eDfQ/AZ8ID5Qi4oEencPQmlCdt91tXKJRCbH0Bj
Bb060pC3xscFLTne8FHNwyvGYu2/+XrvZVkfa+wrkIkLugBb+jeNGK0SOC+DQ6h/05RjTjqKPlcr
hAMblZCoslFM2Zzt0rT+/iwrtdoiAtx0zDvsIbOMoogi18ZBmyZIy1JyJh9/e2WKmf5PUq8/sWEo
usunT+nas2iYDE70x1Kg1dl740HSxu8uMeCOR3tWduaxM1aHr8h4Tva8TcYHMQFFLUbpwOk4aWy9
ChaI0Qtfi9VM4JPG/re55nOtzHhnu9+OhF6gj7n48898yVmrWa/r0sqXP9dHnNCKbVcaGX1kX9NE
ZCWhvQefU+iz1bfi+hynT9Iz0lXLMQiUe7kIjMYSNF9vvPFq3jnlaZCOWsJnXUd3Zkq27p2nurIp
VyoCTUqxPLTA6OtZK/A/HmirQs+RS5TWPITgCHtwKhpsGMysgD5rPV1Vl3igE1bsf2EzJB1EUxDs
8p1634jMExXazxOztro+ibi7TFhmIecNeQNjdLJqI96Eb4d0/vVZzWZuTXIPjdq2zvcSiOK8vJqN
UBsFsHjf0vVW1ru2g5XCojPFvei7zN2xGtzOEErYxXdR7XgtgNw2Go+LX523GuZ1Ve7WNe/rTLmn
IigkhMNCPv1JujKO2XARlGJossJWdo9zmGYWt24m74OqhDwJ6xxMW55pwDWAG8nc5GDKvFtnBc50
JQE4BHpKoeganpUUf6+MKAcWoizGvsS9epdZ0dDn0TxlXD8xR55UcYZrt8147LsQq/FvHnmltK1V
gUgDU9C+QCi6P10T8D1EAKz3HPfa4u/uNNqI67+zJDfr4oUD6to/GjLE7W7Kd5cqmgQP99TZyNC9
yv40AObrge4E7i+JaFgc6tSgxKu+WpqSWlIIBpnhclnKEglGeEn1clB5J7/h4tpEqhsEuY2Elenx
9FID0sRcdbFPFTMZurDD8EYeMTgJ4KLCH/p2J8q6qbkYQVRE7kLTuoWvEjkiefwy2U/GpAVVC4Q+
SwOKt56KTwUGkYez6LPQD4EQdzpG0FnvaDjINi8jL/aOk1C1p0QlQKqg/z1lcAOLIBlIZY41wrfz
tTUq5bWAYM3GCi/fhcW6D7t1V7ChEjxvpColWFvdifKaeCNQeiHQ/BwpE07WPWClPKVm3q2X35gN
d8amJUr1cJqfFMF4RZhiIeU5Yvz888Cl6MwEpZnvOzzwvZxv/yOUVCPHaPmsiKo9GNrq5bafAM4o
619wRBpMT/5NMtzTV3NtBezwNe5ZFMxRv61GVPjIx9De0clHfoX9ggjCAFl4gfO65L2xHcu8EDoN
iRS624XoCVKAtFnNlEhXko+YGHFRBs+EQM5E8wEHHbatcZIi0IAmuiqsp78NHLz9ghzT2mEp1G/d
tKX13VPIDqJzq+NhwAvdoLEz6vnqgB0FKhJozMiNoHdwrum3e0oBkFwuocHr5LXFIhPdOhdAYYsW
lftvFJkAaRQNpjoo9ZLGtPMUEWm7fYBOgJRFjeJk7U9twj1RXU05n60rLWSnrx4sc1L6b0cjHtCx
+hIVvUhUy7Z/jwI9a6r4/Rj8MSYVsVhIsX8PxISl0fhQZsaisv7Ca9WmUkas0p5kVeT0Caljn6AX
JLQfmwiSqgehIEoZKN7taIIrn4W8ERdIhtyYNUjdpSq/DtUsqxX/AgY66QBLH9Aq5MdXWdtBhWYE
CwcHl5NfM/9apzW4F/esqj1kUBXhcPa9Wx2kcrY3r4zcGrRv2JezOPNvySxVr074tYgUP3W4TYQe
THmXSSL3vULtIouTF2swP3rafpt4y9Dvb4il+LBuTu09rKNbSo3wUgAgwKk2HckPyjgRI+ApaxGs
JTlB1YgHS3X5tZ0fmEiqOFMVaDSH0mTCyXevAUKsHxUia/+M6yuFNvTIZl+SjmqnIVVBpnlU+wgl
uZzH2NALs6vLngq5gklmXtQK+/Vyx5/KMhaq+QHfdqV3sWTohxbf7/vgiS+gGwYnQamI+DzGU6KN
Q5FjNZzpnN/7wtokI/bLuZgZm47y0Rkqy6/WQlaEMyG4qpwDU29MUVPA63du/sGB2Su0q/1We/P7
QRPt60z0K43CyxLgthK5tPdrr1RwCxebAksOLqcCOPCnSIecF8vimxVuuj+9enEe3s1F/dTV8l9+
fN0w6rN1PG8fCxF+pmbi+K8iFTaaruKLdbSeY5Oy/vj25ZIQA5aUUY+W4YACvAKwf6JkPETdOsXT
Tf9bxRP2ot0iMBJmfaWl+fnd7z8RwszoJW/2PkIk1bt3ckL5/jA/9JdOI6uE8EM7DcQ2BEuSpnCo
qd9M1wdL4JnOf5F0O5Qb9FFbPEJLKYI1eHJBpWxyObcmFJu5MCKjYv2ooshWx9TDIdHiJHTTn8Uj
RguYX8VDtWimaPY+zQBzUfo8LDOB6oXJz18ksp0euKUzRuMZGuVwBFLpeeekphtzKneerJNVYKnb
kjuBdubgT2HW6LlPPXa3l9z0nWb30SE3k4aWe5QqdpKXCZFHUS2/MbQUcTnI60T/m//iq0VmOiLz
ZyGEamA/64aqHDTMdCCyywMBrabEM1jJtIFOwCdakzcEeWIXHwj5zIW4jYJKsj6FAjhFynF/oITO
rgxtuOAhNtkRDKhjWVa6FwfQ4mmItjpsa2wUktdiGFLP3R/nnutMLxD3eTfSTsFIeKK+4e6M2Z4M
1Utm6Vq7iuyw3xbyZwD851q1nG6sbAJoYkygsDyuPEOFpsjL0FFjyalYMAX+5r2Jj9oo2d8660Bj
G0nqmLlGWLG04uOGgPGOoXPYbGUdgo9aHBzd3+NcTz5hp0ADSENpQolLe/FKACR7k1jd7MG+6IUk
LxV076P7K4mGbmP9KwhAX4HPfzk3O6TXlVKYMicudH+bN1KG1OvV3Qor0AvBbh/bt9ndHmpOkEqE
RO9oQQJSJwLxB2lLqP2OyRDJ7RyLW09nujb0Nf32WikMVjaCTqTbKmSNLIIkqDRXbt0E4W7sbNH5
0VHqyIRDz5253D3UoiQ2oI0Fa1puc8B1rDaahsTICtSJOyphqtpRzmNTdBdRmGw2ZNdesat5PHI7
N9BeVJcuIhg4pV61v8gwIQGg+qhSkpciHiz/hYDv2VdEWveYomLLG6R79y51xkLMnQBwBvGRSjwO
HWEgLLMj8hjUKec2ONsxALZlPk7MCMvyDam+87U9m32Ka189LDlL0D1VRRim5fJsRey5uPSaueiK
mBfhdCPdLffBYwmDjZs7VJWlef65LXOK5o3CcaL483HVPGiRQOY/BZEmi96E0SgQJ/Or71PEivs1
lmLzxCONeMORywWu2Rv8LXfQdFi6tn+hDQLLAkyLF2xO5IsCpY4AzNDwWoK0XrH1vRreHYZCa8Fb
68azQV0nC7CCOWgmITFbs85gv8/FoevdNh5tzJJmfHRpF4Z3TwfrUf+UxFJEHXZfR8SFb/UfJJOS
uCyt7kUxbTxC99KDYiTTQxWKaqFV/ZWc1BD5ZtXyn6tDZQYfWuF4L/qyzW/Dp0XuQojCyRLi20Hy
TcguOBtar5ods6eTAziqz1bmSGL8hrGHP+4SF4Wh2kskI5pGu/cI+eInqCSVCI7nIMhgU8hCNj1U
zm8+ffVAnB1/CJVmTMqPEFHUw1Qv6U/2Q9R2JDo1fB5h/HmhVZ/i4IKQZvwqlIZOO2fZjOXyDa6+
Lf2SqeIddL249NX4Nds9r805SjnFOdOQncSgtRBAU51CDwTCl9iXZyRVmRl6hxsopX+g0fCWVd3t
ZZlqTE4By52w3osPXhkKPTmOjp6XEiL6BgE3qHQ9V8NJKTOyTV10wQR0MR7Qmvzx3R7WsszfZDw8
34YAUjm2fhcwMptsKu/DVphc1JOs9e3OmSRyRktybZmPNcikaxRW1sBMYLkGptVYsFkXX2Ycfd44
Y5rOVSWgO8v/S9jfBUIOF6E8aAlZ8rRK3StChzOtql6xwDzhUyzx6ivDVHEUSeIZin07AbnJPkbG
1eS15sSbM6sRmCYthxGHiXZ1rQBQS4/0C82TlPbK4s4BEmCZX5zX3jbYUA3VjZhdBb0hiSLStNTc
RxSg0IPOCMZFbnz8RmaZU2CjtV24yl9GWRdxs4SskxOSLjai64/MYg9lMWAlMoXrVKHy0nJCFsIl
9UpcXq0JkWEDoe9iQvOyTVWPKs8BcBeqqnh+sGOIn5282bGKzVhdL3oMRGH+s0HhLlTrlLVNhgkr
p02XZxlvgkg1R5Jo5KDbjz6W2+EvZweiF1Ba/Knonbs94tpxOFuXfK17zcViU3OBSj+8EIfJ8C20
mA9nYkqyKa4c4CskplftJowxRP7rRhFsqRNAGrVOxV4WS48vLedAjJFpev+2jaxCY9NmgdliTkqy
wpStAtYRIpK2W2kGYmjvxu2RP9VnuEwx/ANXA02Y7nltkg8Uv5FLtHP3Znf9D6MTIJmO3q5goL38
fvx9/qxUxda7ycU4cD2nFRiL/zgUlVP4zLme7pcjbF1dnImId8hwx6GxVEoF8dind37QHpdHoPNk
kZT6Bm3gniHUaHQYQYWoPxazsEXCXncw+U+zkK6V99y3I1CSvMXQQFCMJHiIxFfxnn0PNyRUO3OT
moVvfTjgaNtU0XvH5K+UWuqJlJtslC39WC/q/yEU931A2YFTY2plCVmoTlkDWEOSzokSmknZZwHe
IdFtn2ICKN6wNcDLe0fDIemQ5L83VRCFblgQJRx8lJxa/H0nLCQjUOMap5+zR4Cd6cAQw0oZQg1s
4fhvXpCqEwrW+2Ncv6FMyxOuFo8Z7jpajFtLLGO/ljVEO1WlBtAfOGRVWyfBn+htvW96r4cKtOyu
9e9uctQxybDVjExHH0T/QbJ2CNSG/m+C/O0R8bB3wpduSbLofVyQb4BpfcRoXz3Dtifz9YA5y3/u
VnZFiL8qxceJhSVXMWxPhouEgE0qMpDTOCQAcMejtLzN9rXLEWeRvmVkWU/IMyeDKPCFm2fbB5d6
jV+D5kUaqvu1aahetsrnjnD+lP9S5FUM/bniKVzEmOqG63DezpOqly4aFXtgvnBc38q8ibtLuaBH
lcjwWPMo/3YJqaiOVYV/jWOJEgW/sM7+rKlWl2xcRraur4+Bcp5949DQ69EVQ8Mvxg7S/iBwNnZJ
FZtt6yMlRe8gMLFCIHg+E3TooDHFhowHF8djRvSowHvbQPih//67ccb0AwKpKwnR2mv/iBMXgjv8
wm1JjF54z4JDCVJ+H1NykfcILK1lsnOGGtfdZ2Z20PPXLHoA7oYr081ZOhXnXKyBFbM0YXLY5moP
WJ5deND767HO6wMRoaXpHIP2s0jAi3FHeQ3hYW465GMWxMcECeVJ2iMYVnTa1z0YlxYwW2i/DQdE
qM3Xj7FiilUmDO2bCi85BsYJcpBFZho6P61LnXkcti4y0VDDEprcIZJIml2BUDsH3OqoNhyFd5be
xvN+3KkjIPoAHwR8/LSnwUaIV+K38NlWW9U2ZnaK4+5tegc0UcI7EAkl8oWSr/i/nnbe99jUJUkh
ZbIq2goK7mcD27OaaNfHSyXWyYhKP3RoRdIknzR0G5yrUCLgva8BQN2qsus5Ast3e83qzfh0PLaR
ATkYbYK8mf+aQP98wgs1QlQ9pjdOFFRBsNscqaB6I/DIpA7UGyasshv6HV18nv+5XltxIf+6DZc3
Is7of+hblocuvVQiao1JnKNWyLahZhJt8pv8VGSXxYxC1GUW+j7DCS7M5KMboxaB6iE9wYTtEpSK
glG/flv4tjjytWcrD3EdvyVmS1OXSdFwvpun890XAnIwQYJMDfAqbAFwkcd9NtIOTOpb+6Z+MLud
LBukQZPNFS9ttVtLRZ/1uVkQAb2NuLU3zXZz6NcZSnqA1d9IzsAMARQN0sBkbAtTWZ7WuRYrfbYy
vp10yUdpLFnQ/z94MqP8hLdFFMqtHdu3+0s7cZoNFb0kiZOp8I5rgsjWfs3DVivjBTu9jkmrPvlH
Cc/FABwJrtZ6Hlo49U3UJyeWmfitI+gw6UJLR1rpc5zy4j8ZVBITBKKogo3Fylq92Pw3BW6pOkYr
SoH9IKu2mbq2vJ0s9jTv1ihoKnelaYYmE5Fu6UznBx/O/JV/yM0He4tSOHEPztYgUzCPiuIpaxBv
b7s/75/rb9sI03QsOBcn9uFxBzJrlCPHmNQ3zLupTYMjWyFqDTisJVqABd5BTcB1J4ovgjHJ0dzb
gc/TBtgVY020NQOjJu6NHnnIQQCNa7t+9blqJEgRNCqq+FsqpV3K7aSvKFbrfdrnAxUqnFpZumN/
HEQgalm+XyRohhdFvTSw26cdbqxdiv0QUFR9qbBWOYlU4ai46M8NGrvwvgBDV3/anhQpEBG6b13A
IYaV/pWkcc0DLaPJmz6abrPydmrD5Fjl83uh6bGnFFhLSUrPmqmSiEeaEogZr5xytArbb82x8K/l
KOd1blIOC7xm08xgNXtKqL5kH2BrsCBzfx4fdBvyR90H9VA7xQAyJCOroLBooRCQ7USj/mzR1NR5
9kIW8d+hirnBWeiZ7Aws+DVDRsGPBVa/oTKuLr1lXefa4mdpkH8D+UpiIDFD40NiMtGcjTr4eKvw
RPk7ohP8yLgGwUVLdFgPssiUOS29W3LYMPq/0mxRtVxmDM63T1KNx99ypGwmU9Kx0vgTyDVkxG6g
1BOfam57/Cu8m0PSzG7XOtlkNb4y/vthiIzVkTkWBPsKGH1qdwutbChg8qfTEX23D7SXzukXs0tt
2/bIL6c8EU411mANoGLlG4132Ql9HEEy2Q/M60OysVt7M4JRBP7kZCGvAVAT+apvkYs2VUtwPWx4
Sg2IJMMq76zRiHJ4w3WolSurAfz2AsRvnLbJI9jq2am0S1DJ2LW6Nh1cOS1gzi8LBwEihIBKilN0
6kkvz0fg2+QJkmEAdnxusK+OrPyuS+sFStJT3J3+p+n/pzNhp0tignT+naAbfD+pe+I5RF+cby7r
uRgN+cUfI06kpRUqybqgr6HhxVr4gH38pPSCJR1CzLqAIBbJDEfsafbDXhvzEOill2x19gqu7sxi
0PLrUwksZQTHehBB4BNNBxdiIDdF6GHOWE/qAcxxPFqqf31nSCpe1cJ4s5AHv+ODiphTqpK4tmTK
RSQHR6K76ntLyI9kWTeM2T6Y7TmcNS0CkEP4KNFuS0aKWxr+M35mNsvjzbFqtp/WIwtS873k7CWl
X5ZTm9Dgs5XSQSGZoNGok6z3cWLj0ZbupVK9Rtbcm78qBbzjibI7xGn+E9qjWEtm2BH8g5ilZuY7
q0XxNbs+nAZ/pZNeIOmNsLPAf1f+hpIYlsTtkB85xWBkEYmRZqBsTymSANpfBHptb27tyS7TXg3B
N6RBcMNe50ZMLhNGiQXNbxi+iYRpWX6fHJ9cL9tpBypBgVOquU57D8esRvchJAw5gCOVUiZ56Guc
+vwAaTQSx1MIxAcmNcuQbxVCluw6sEKiiGGCz/G5ficlByrELXij68sHnyuQW0Fwzn5g77mkXIIC
igd9v3GPxTEmrsOA9kyN1GqhxGBIvjhe9VB/IWGvxtnwXOrh/Q+G+Cak+8tVhmxWYpYDjL+4K5Tt
eo67kSDKWkO2JBcoAerkRYH2Cw6DHTCn1YlcLQtNRafmLZo/XVNKlUEdOZN7PVncmskbISWngl4n
mbhGM+OgXKhayr2ssB/VWpY6dmJKuTbCZDZGi9htVai9gjE3Tknrfd0nhfS4yvVgBhko743DQQ+F
rgvuAlPRhuqKa+umjIPBJrX3g+tc/FJoZCpCrhzmsV88woNzyjEVjYKejy42TvBO1azWEstWY6MV
/Tj5Ofkf9wpnovZMJonYkS1EublNfTQw1umfHyh61GCsXawxL8SsKYrx1fsC0SmQS0nO1nsj/zDt
H6lc/c4lSU635YRqnMM/0Ss2ct91H/QBWU6+qYBH5aue6/P+5GZfASPgJMztLutfDrv7aTxTSYaZ
+JR7dlQ7b4u2iAYdV+CnX9o64R+eZ4+ad4dUWiVs2vYKYK2ySdVReIvOlHvURmk214a3i7WUHPO9
UGlndXms7FyGelPKMGJRZ0sVDxspxirOiWJTtOsROd0ViuCY05ESIjgQbD7XyW7a56gUzJ5c1/dA
A1Znib3adKAihDONOn1innuGbEX112oJnUZ3mKMNQgUKIG5c2H9ANCSuAt015ZVQoGFNs8TWxffW
sEksqcu3Wyot87Di8HyUGvfFGBmzP2wF1zDKXl9QIzy8wdk10PKLmakpD5y3ws2n+SMHOINwzVuM
Y2yKTUcuFEOBfDUrgVPX3sezUEiK4nzIR2YY5RDC51Bo9zNq8GgDIasR1MVQmeCR7R/xwX/VEpH9
dQMfEWE+pbvkRXCxRlIgJl0whvO1p1q8N7GKmvMOnuzQhcXreMRTQK0DQDbx/6Qff7b6AQfAeSB1
vkcmB+A+3Q+JpHijO1WajSKPZ1zqKOKexZdzXLhiTBXUj9DnTjD9QMTZb8ity89c5ygjBuK8kDEx
w2HwHouQy4Ztxo43iXQ2/oGbcrSslnYfkBattUS+y6nXcgvSamr+m1AEQSb+4WBK+fAlrk14UYjJ
0a3tW/KSQVxuYM5Me04MhOejCQ/VSC1LNJgSc2yfMm/kEmqsMPekiPPKy0V1J6HM1djjbTnNDBiV
02xkw38qdD11APlPRpAy5JbGDqMp2TkieHo4iAQAJ4/7e80V93x3jGtjUEpVJu0LFhoE8XQwqstW
kRQrZlD3Wqfi4tej97tL7TX3KbkKGYiTwQxoQfAYTCuzkl6YmCb4JS6x333ZGD+TmrkZH4jX2EbQ
PS710Nmk66N2j+9gyezRM50xfH528AqXEdz6k+4pUahyPcsr1Z6G5d5lXX4NeCZdejTtM9/aBTyD
A+jM31EOdS1NzHZFUIFhB2wPoAc/V2SvtpMZwpXLCNftKBwuuZp7SIU/UzAvo3QlDcKuANKnN3Ww
htlmS04gDdDxnrb4Rct4dzSDGd5G8pIbkaa4zYBT3B1RlUsoyWWO14AZtXpEEK2l/WszdaFa85c3
m4OlfYNHrexSR4lVvukGnW4V1vBinuLyY4x0BFYt7GEUNJ7SsSVzLA52ru9ugseWDZ1uP1Gnzv48
qeNu9ENFIHWRhzho9b6CY9bDovDeQ5MDK3vxnLs6Ek+uOMUNttwL8bMtIO6KbR5g3wPo7GQa4q7E
iCPzVbVbXI4PDM7SXArN1qWcF8XxrfgZgv9B8HI4c1yZR7UzUo0RbI20RXvex5ii1JQjPmwCx/1v
B3V6bvYS5XBj8BKSiwp2rBcRAA1mI3jI2bJFzGx1Pc9VfPRu9QpuEU/X+2GjMLgEFHo1NPuobd/R
eJbtLHEmSjZNMLApdYi8MTP1FpoO4GoqRGvkgpdde1jV1meCiEV5tIG2KjUgn1px6PsdPcPDfSu/
jlL7lNwpbi+O6YIBbhtHR4AVE03qxHY8vX4D1CeOE8L4VHvrgXz3JcfX11hH/ABw/HrmTIa8ow0H
VqWFo4Xq+Cm7IIm/k/M0bLONVXbC/tp1DdHh6YKX3ZmBEg5MeX1UneT6glj99sGSe4gtg/jHtTvt
v/eE4TyTD8I7QopYvNZixG5w9uRsjY+gzSSJ6qgXdDDx+1DVdgNqY0N3EXJoJ/L4lVyZf6f0yj23
+BjOsi0FC/gb+W6lAdYaEEW8QvGpL3TXYvDx67keItjD1K863eiFhV/8rJ44kN1biYkExJ/7i0tJ
dpWEKRS+Be623zcO3vcyCeMaUO0KCv0gCl6OEx5Le88M9xpIeJlpsjyFVzcITdo38gs6xWedzZ85
UfYJvbcQX+8GbJasbc/zHgsjW/qLv8vjn+udilF1N+uKuOZVRhbLHV+m5kTYEnOgBfSCwYFUGhPv
cFRQBLGlYYMwmtiPy7HKR79r0xfYVWqTMkym0SZOCaMDSfpbm0vWPp4ln1nby+CPpy9aqyekqalE
jEqLoAiPMKAt6j94S+s3qXZ94Rr4Mpfxt+gddkVfuxiQfXM0sRn1ZtZkZxcWUyTVo1p81bQH4+Ac
SjoebRLWmydeJMoX4iqQLQ2FX18ONzEwzJo0Zsd0c8hNSO+jeeJEnrdNLl/qN+NrMKE19J5Wzw2R
RGe6uxK0QGJFt4exsEWS66a1Cs6ZALkxgYW6EFJhhqPldZ18QDtIwIVWL57kI/sN9Hb1+5d+hAIE
Mibc7H3XGNJC1BBmlKt2jS7u883ugdAEv5Y4T25qx0ojIxTfR8qcD0oYG8Q2uPP6My+TMU9JyDUp
M3GnZSoAoLMqDaDC8VoOzQHoHS9xv12vye1wXngMwuyUCrXx4q7vWZgVEAP5S+0jFzMXOxOouG12
G8/HXKYyvd+gYwW/VDEwgrdrnzfGJ1CoJ4ShtPhr5MD6HRpp/qNEqw4TsrgS07MqCWwDYL4JVQQi
1vOu9HSKGf7d0Qqv2FT5+ozPq582fRLAb50qPErQinMIgFUzThRgRrFT0wQ6NxmPHdb020eH2SCg
wOdMy8fct2DntttNrRMnP8c1G/nILLhZU+uYmMJGVPkyfmg12bFDn9R3unfFZKxexQf4zh/78UVn
SDtE2J0P5POfV5+qD+kIQwYw/f+jXXVta/zftNxHU88jxzqASbZG+/ZdVsPFaH1QgOrizNqtDUHB
apC/+8vEjBYRWvAu8yiD7Tus0OWFPbREdJnoYhjojkt3SIt8jpMykHRuaCyt+nFx5j+k3E2vMZLY
/4Sk1mAP5Rsb9LcL+vMlUYPIEKe5E94Qbc2yr/G7l6+FRq91eBU+WjkguHEhWuXs73gSwpwMpC34
0hguV/dLNrByykhk2OMMuAPGD0a1zaGgWp27iRvwry7OK+Gig2pkFuSOH6SLkJJm25yiUv7E2Fvs
jnrTmy+N8wLaXJDcHr9w/J7dP2m18kDwfrfMgTuwI9ztx8DpOcoY3jR9wgYKTmxu68xl6FO+5tkW
xWdB1LryLE+o/HbduRYhcyVdrPFxDLKj8cnv9CNpRXfiQY8UVRxewbhyz+WLjyBlBqnj3HwuDBR2
WEouOanHn+N+2G8v1EODQDAeLadrh0S4hRQve1+m6yTPNV/RPfpPo0Eam498UkDXJ1K3HLRYAdLc
WUV63O6l36Jxaq6+WABPi8iI6t5WDbI+YTrvhVtP69kg0WRaNMVwJ2dy//1dI16ywB6JKUimWQNJ
ZiU5ZbWpMF1HgmLrRXY++MU2RbWZmmdJG3xc7P+i3G+MmmZxV7pKMSWi9lsSOGkeNf7XdEV5Km8n
+dzwHKxo5LotaYKMn+2VzNTD2f9ATKbBQz2rzx4mVUn5glSGW1s8+dVeXEGm0Q6qR2y7JVOybq5x
F/1Y7LyXldvbP1rm6o9PL+qrj3DQnq8MGGuXr3metpI4mAB3aujrQZUKCauALjTGQbiXpJH5rYpH
ULa+axmCQ37xV+c2Xb1mlSgGXMNCL0FxEtaXdSt53RUiqdHF56+nIP3VcA1Myyx4ONva6ourD/Ol
6NA3ZdyXZnT1FuuQt8eJSbUV3io/9+v0TowHQ3Q+cweXu0MTuLc0N3X5gv9JNeBv20rHieTZj3iG
khQ0AIHMtReKSzqK4Zajam9M9dwqjI0rJ54iwe0qulegDakrR0iuiPe8bhZcjl45YyBrm3+X+M6V
6EzpXTzBXQM7KqmgzHSYbVYz+o2A+TIO9Z8hGoIJ1h/QxXfTuqTr0Q1j2ye8NJLJaqo8YPj6sKjk
q9bsOkauDc4MoO1dJkeRjROnhYY6eaxCeu3uh/LBCOHRKJK5/oroEtP8CfEPVibvtUM0Z3ETrbfu
fDCNxK6XrulfpGhV6qRjJfxC/i8hq5T+YJYN9Vg8YFMF1Uolup9PzK+2pIGQDh+PAmBhe41MIdv2
B8nBLq+t4Vxry2rTEToit27LmEdQ6+V3ZfIMhJ1rkzh6gZmsYUh64eI4tuwHRR+BM9C4R5s+mIKH
+buZnN6VuVkWS4l3UMlGePUJ7t5ExFAjp7nbaZDRWv2F7rPaaAxhzfvz11t6KedGzBfrrQ68h2J7
S7fpEfJ7AH4d0bnU9uGU80qHjyaSqymPLKNbua5QJkG1f8cTS3h4BBq8zL7XlHL2KlDm3f2XeMom
x+FW6nAD92UDDuyMjk13fN1KbeYZ/n5Q3aAooYVad+3RbGmZ/oO/jSy90BWI+Ney5QYh8QT6j3sF
5J3CgIUZg4o9X6YoSf+qN3X6E0ZuRi+20GmVmHW2vFba6dVNfW+V+eFeg2nomPKT4kGYZT0S0OAK
oPgk67ZGQXY4ilAVJDJmSVqvVQTl+jFbDDLEQ9HfBRozsflaP57Vkd8zV88OhMQQHru0Xottt+1j
hmIh4c+92lwO3thyRVvaz6rLWyPrmehHWiqCnoaHRYBtXarBoJg1DgFZp1Za0IzpNjOsCWFgeEK6
2LZxAmcmIK87NM9aEis16lTdhnNVaJl7/jYjjbuDPlHmfnjq93XK14nViR8l+0JFoRJHJyStchAo
hgniT2mQbC7DPDki4Uec7kbKl+vqwTDyQ/uwxmPubKzo0kUI025uPZo19f9KcjFUMA2ygzN4AYon
PH7eKWgGkk8Vc2GqvJzEzrgB69gawQLYGeeGevvttfUYfXq2zcaqH/KlXobmsWlAw/OpzgmffBCc
qBBK+XCpBarcjLlynkSXk5QwEV21bbYhLnzd3T0vg3Lw7V3Uhox+fPFaxeXsKesZ3b9PACiZhiiq
VGyEM76kjrJ1p5Xu4NOJb5HD3lK+8KGhlVuVsuq7DoFe1fC5aQfNWvx+If7dUcNe3cwqM3Z7SVo7
R6Z6+rp5tbAAlxRIbD34ofRxo+FE2tPJalU517ubZcrPNCYJkbxOV+dTycaozZAaO+pM91FHsssA
Q1AC5gqz5aFTyeMFsgIC/qHwWOyjTCQCoNxs37ujDOR9jRjZ0atKYPGX2pW/n8GhUAV8iPA8oII1
vPc7WattX8NJlGXOMmFigQYViBWXKGg8AuNrUPZfU9Bgfr9k755TbXTVh3wYCY9N8A4KnOLr6X1s
+0WdS7YccA0qViAqviZetT7sfAt3YJzeD9FCcSsdGhpN8LTLuFXCHurXgOz0dVvlaiD53YQh4OGs
SXzBMUZFIDMfZjo6+j0f/MRFa6d8WciEn+Me0oOzae4BjkS6aYyUlJriKjQyyuHlZLfY/5AfMUYD
nCcBHw1B+y647WS5EUHZZgCr43ZsP0Wk/xTWxeXmg8RgAoppHFQ3/XFLrGn13aPwbwf8bSfzE4jS
yRzwrOl2+J7x6mNn3okO2K9NjkbgPDeM65TpgfBbRjJLCBOw8Lt2/47Ukm7V8+ccMERrq+HX9wx8
c04zs6QgwHs+M/60IvaksRLKzI0oCnK0BL/MDla+45QFCHOuS+t6EoWZU7/0J3C7YOyBW5xRaei0
Hw4VcaBU5HchO2t2k0jQbgigSdNvPZjfHxpoGaFi8fQPiIYXWII5taav7Cu40WWVCG0jjGPIM0Ls
Mf/590xX/F0Mfjchf5geSvuGY2Lixw1J5Z5jvMPTn/IifDn1Nb/yf5UOURM3c69K2TL3v6TEW9E8
aTER94koQxhgciJ4QXtSpy3L7/H4ioKhc3ktzgeQgfR3AFMsCpN4SlWNyypkk+cN/WUSlz+IKf+K
J/K5Hf21VNpTiD+QjSDHDse0oCefJLuYHl1K35EjwBKMgFt6fwG+pZ1NjoXxdDcW7cA3rGkWLwyg
8R5v6aqO2H7zz2i+M3IC2GC0+fXg4Dz8b7yZ1vRqpZaFzZHyn5uWd0Ltj9SDcvl/zWz5/x4tCwK8
aLkp43e59ZfC/t380zInb/9v+x9wUctgFFpmAguXK4l1NT85Lbqs1a6ntMuVx3tRvyrs3oPGAy/H
ke6r+SQUMTp6OBMAbZ+/eOZ0ZDZgtJM1pBYNfyUbIBRLnNtqXTZLaJFh/LFf8ZUVKc71PF3caSHl
WDMn/AxXwBAWDP9v8N6DkIPgTNVe6ZzTAqUr/qhqujKztiwIOHR+YmSs8YXDtiIk7VTYi7oWUOMe
O3Swr4VE7DfsHxez4TWdA1cCAgAUYWIOMXBA+yGRf70DZUpowD+9qDV7dr+9C1sku2YbviH23yVA
cSS8Cg5YRgfGItjkMk/VsG5OufI5CbU2f3Ry7CtABvcrsz5nEI5RDCQYwZT+nKlJ9AkcEaovGEeb
DiUyWY8FcCOOwmzhRINeI4uoe7dmPMIZ+rlP2c7Etv80tfPLXbWAFnkf/MTSG2+giesXQ65LL5vU
1nh2jtfFwbBDDuNvvRLXg/tEwIAnqw0cE3EMWSr6YNceOFcQuWSJmWREERqvNh7WRqiLmkoNJ/Yy
gWDwxvCTscOiBxchdh+Bfin4loeOrn5+jAHurQKLN/F8cY5biFeFzFXGD35fKWljYyh8ik9wDIvE
buFovwUTw4a5FaBI/mdM+uHCiV6Uw8JPF/9LmjYfKrkO5Wb+2a3IF56GFhJAXFruvjvGbRdcCtM/
8GwHhNCdftRXD0s2+JFcgbry60x4pZlVGyDcWUNQ8yFkNXFyvbKCu2fQ6kRt367H+XKublFUOF3Y
HVA1Ststv8rnlqVDpEiKgDpLxi1Rj6eaRVYe+/3efYsaObiTQmBcCUnvGa4VgAvJ+OsHa5EojLVy
CYByy6ybE07uU0IJY5GmTr1/dt/UFNEJjQLrbiIKjcLOkTO+/0RpVHWRSg3Tw7xvwupw2rGkrio3
SVq6ZhCLrTcb3lf9ciW0JZuHfNr3S+HOxy1FKQjOzzMSpF9CCWQtztI7DEvPSaf0EHfyseQw6ity
RoFCXywwAR6Pl6NNQZzVuDF1InqSIXgy13hlzApBKRFUkeE2XcXfWwbmZ4a5OM2GjBqXZSf2biC9
Is7FqYzWl0N6GZSUJtn5WySfOqUn0FKl+8dZ/hu+YiP4tgqGNVWPYvX7edBgOgKJ1ttKvWwPhY5t
d3ora0UfT5NZ/hEZauTRvpiSL2f3VI2Kz+mJCLPJRey7mgTwYBgJotUXrOd2uXTZpLToN/AW0O+V
/gZAwA4GF1HSPjLwwE1MwJrJDkv/AZlOEYtjxFe/87IfFyaPTAiT21BjyNIRldSOUq6X9Sc0CoAF
odyk99R95trh9BwgAACS+gdoFgGT1RQGS5D5nrHc3AaBY+lPPrxMpx86EQgz5xYcEOpiDC5QVo9Y
vtfMx8jNh9NlT83llx0y6eTvjDNHsnJzEFIK5+MtZIhLHgjNixCQxY4jjh9yHOa3uclqMwle1GgW
XYrvp5eY4VE64jFJkp1XhMCNqZLVZi7GXFpJqjowtUIkgCpPa513XYomhL9dC/4f/0CcbpyiFYGV
UEGZCyRz9MVuBX7rwdTLVmNZRMYyT2wcTzeY/hi5XTwzGOjaOI5LllULApTinogYCL+LQkxFhfcZ
/8XW7OmN5GDV7TT5hlejuWnB+7DDMmz0HS1cx7UHJMFi8U3GLauyHzt9kw+r5TzKvZPdVCLlYE/m
7U1Y2TCizhnv+E00mOHfQHbl+08sE3rG2uO91rAlj34L7h7Dc3niDCv8OxBe2YPKNS61DIXCXN9u
nCJbhcB7HbAj8tcCNWq4ChjTWHlnxm6qsuDI84Yug4Nghbhf2TIe42tRO+gB81IhU7zfPBbUYEJd
u4Rm6tDlsyZ9tEvbOxOuDMmWB5pz7aCdAA3iA1XqI8atHXFGiF/PkqCe0HFjB7phTjzY7oCsitdh
m2UPGLoPXNi+m3gQQkPxzInWWMm+N51Lp8yftPrUG6rBh7khKtvg+AU/Ci7W1Esa+qRWAMgVAuc1
BZdPs9yizMI+7ZgrP/iE9agPDHJcEXN1rCXWxNQ2Z0z92IXG96SwiWqpjUr9U6T/dDtF0F+xpLBE
/dqvI2HkjDqghej9P1q9Kv2Uwz3cw3VX4u1eg+EAwihz/23wekcEM6dgvkcu+xTV3bopauIF7/JY
t4oCp2rluMIIyXWnOdfJ5tiGURod9LOHBUogaYkeKFsz2EX5gOnzeTK9VNBhRl65/7qkddOUjvS1
AfxcybfNuzmv9AfGLM+9yJy1VMukBbDtFArINlT2as0L+x9qZDzDRjqtj97VdG1nsowihttu2Mbc
lPhSYGf1RMmX0RbUAW5r6I5WLtfd5VskM2bArQjmwvFy3Vk8M+hdDYInSPif6Y1NdD/+w4gIaZww
vDjtT++0B/MRqNt0WR6E6Pm4rABaBiQraaZcPG3G1/4RiNZot2g6KboBS+1d29M1p/1uJOTHHkkP
jtbhPxMZfXYbGyYMq3Vp8Qulnly5hVR/5KlOkZniZEXutfm5Nkje4uEPnTlkHljU5xSRpr4AMqTY
PeMpgg+lJqjEjvflOt+y7kEVAqA9bbamjdK7FBagIkAVvO4FGGH7iqPA0mLgnQ6EOVvhNwKjOcSa
aNPEc9fHe0E2UizGVIKDObLHh5uMWuHDeZDVcJdLw6fxyzBhLqkU91FJ+z2qpANkxgptZ06esNXb
RgbyICavwH+B77kMndj2+96OblFS/2F7Ge3X3fGYlseQsVsrCjEJSP7ATxSabRVBhffltrHOKdbt
6hw9IGcr2dQq9Re7KhM45PyBnJt40PJLsQEVxwV6PsP1weCQDJP005UzXx6q665PrBJc/HUTnWKs
QQFKQS6gwYnHGzk35Lw8LQV3b8SfoIQ1T/KIQAvxTxT47kyUwhdZFi7jDu7SeSXurVL/E4OTf6YX
6RFQp+Q4PPhv9/pFFLI+0LbBzSwJJabkOJSQe3ImgAS30Rwnt6C6B+usCiDu8nQE+JfKjKCtuPHp
4NoWF8lH4iBgpEkkNCPDfmSpnoL3UHyDrWKKQxX6qSqPNdQvxiccM0sJJwfp2BJE3tipWnFreRCZ
99RjlzZjebf/k7GGtyTwsHp5eNCY4r/2B1hsrvgahDlQg0BHZjLpUkse/4RYyFAVZ2kcYxWjduXL
qK9hzzCk77Hqo+hCcIH8vEwBbN/ZxjCYQXKbRZE6bsz4YTNw7S2nmQphi187pJXk06mCm9nXW25J
81ghG6y36/j2133eMXmvhz6ocDK3M3nMGr25Zt1pZ4421ia4IIN5lsVA+gLAKNHg5MU8wr8ahfne
Ue/fLspbOgctFb0FIECYQ+UoEYCK1yEQojFfb11ny1h+FjCsN0k6LnBpXdqb2hENpajT/lJ3Xik1
p5iD9C/7GX2dGzAjpKBa42b1nepg7a6hJtBRMHvKmzrgZTzShx0Apv+ivrtPmAoQGIop7bNM1ZgF
/Ii16fH/unqwWaw1wd/n+ulXrA00sN1f9nb7qenw6LfblUOMpAM2WcFAwEYuk/uUgtPPK/ZmbmXx
pN88LGR+6ticd0PmaQuz0AGM71QSJxxVvVbDCSxZ4gtgvCh8DlhcZDq2StjiE7FKcAmTnwrgUjG1
wg+jvvn4IPoaTHBb5p0ojp7K6kQ72YLE4qV4HPFp2IWyTqDZriwUIuxYyIvR6Olsc3j2PnKUnU7+
19t99E4j3u1Qigyp5VOfPnTgu87Ep3x5Ex6GefhJsT8wKckRzS1La5oG1EYbj041yB2XdALT4wqJ
dOgr2MTgYZsh4YKlhGRJJmqcz7SY0nlyanu7DMtVD3lD08nQn8LgcGPIUHRlGCdXOoS93zSB0y69
Vj84aQS7aiMU8sJHc8xh5g8FCCiSoh/611OWFWVsltT+9+1h23RMFxeVVh+GRH2OdJFDoYElX2Ld
Jn3ldh/9cZhvbZVvcgnTI93r3qJZhZ6YdsU54gH7DRXcnvDApoJvyvNuKjMsubZL7wo3juAFBrPY
1HV1ULPNnHQQ3fbtBpNPKwrG5DP5S7wDRg1HZQLGJp9EZ9hzSZLYyBdxzkgI4eTb41dfVGSovUkx
gCo2eK6t2UCnH5Iw5PlF6RMzk3LimD5n185WnHfMHrzIuLKl0bxgWCiWXgXzf0AgsUJVUDEXkF6x
Gpbt8NGY+KR0CjYRa5IFQ2H0vDOJ0prUopgTXg6mMtgKnGxIvS/RjXqWX7TgIGH19oS+6c4jSOXA
Qp1eocuuxg75PtF4JyCq+oEZE5vL4DbdV1yt7I41WwWKrZXMxFHrbaBKMR6cUmMNHQf00GIA4l9G
I5x3w58SfI5+YcaArpniVCzxjPkG1fsQ0RQuBmNfTGPCv3zokZfv6XvhVQQwQfytwANRvXHMAswJ
uMpXIV4JsNeK2AtAEvZttzgz5iTbbxBw/qggfVOLJoTS3o3/KuodkP/sYXMpd5zjSyXZN2QnU7+z
tqtmF8JEoS8byRcQ99ArOpUbaOPEXLVq3qXv5ORq3nPhBtheHFoOuVPCZ4UPwSjmq/o/W6b0wqef
TsMgxhu5/CS1HKkcyv29yzCypb8/+UndgBAr/VPMUtO5b/8z97GO/5ly0OrayzAPtmoAWTYelGXQ
chdRMnssy+P14nONM872MOBpcLPL28H72Xifzr8Yjo9nTHgEcO4zmeLuwxQUE4208eMWhkyp4cj6
gORUWkX6l765af1s4hl07SZMHi/jm9305wupINa0RMFYFUZ1jGoQ2HOLLTACmGLK2uklo2rAEHcl
ifvz2lm1ywNWyCKXhxDHuX5GoEVRzce1yA50GUaYgxTFaaE1/UkhkkCV55SCbcgNUgjdTfJL429j
fFy1IL0lAZ9FPEaC0kAP35nJGTSbIR6OYX6tnqJU67XQQ2ffnXGldxk35ieKlw1kgOy6i4wND2Un
lvjyGSZCtoPihG3lgDT4bmpbab7PycOXvVrxyVjHNsH1RrgDVYwGRY35EPj+2bje5xnaoYe7CbJR
S0F7VWjV4jTJLCCunQv4ga9inxyL/7aP29XnwZCYujcVbUn8BOZneq7znCo9LXYKGkdaN9hW2iME
8whAEqkCki3qEPyTnOS5TQKXZfkjEIQO5z5qJG/208xBuuNAQZ4T9E1GdWWDKkL/ShDteFONkQBp
2n1Te1mtwrpKe+KHkzXHlcj2NynAm5BTlZnC/eb1P1ZnBOHvUnKM/jaRmlpfey8HwzTDcvM3+AHu
PqucpS2HSjMRrTmNKIbuWptvRoG3hDcRgo9cAgITaZtCZ7UkuZoLqI034akNbnkAa/mKnyVQY2vM
LLPkGdWQugclasqq8f1+Hl/j8KxvXpimZnYVijXDK/uAf+60bEIinmgANdDdXEbyd2UWRnBogT1L
BgTvgS3CI8FlEMyy904Cghgl3dMEQpQYkSUvCXCUXg6INLFaoyF6kSB0OLjwIRtoXqlXRYP2mRJx
3Qa4gqrhxArWm+OA0TK3+3zxvcxPf4jcWdAk+dZiG7MNe5yw84EzIL3qqKTvOOG1M61Yyb9Fmy+V
2ptul3BvbGj7zzzr4wZnTxclAz6uuuax4bDwihvPiNSPKZDNiECljkQj0oSLLK0XOxSUctZ3t2bi
f+iZ3wJGM/wXuH3hYNHInyEvj1rcqE2kre3ILAAPV8Z3X8Ow6X0M/NSAiQQKZ+QZRr/4NRBnc3ZC
cb12Ben1vOB+di7dzpukglyPd3tqoRfpnOfQzW9oMOg/j7xtQM8udKYUiFVV5hCmn0LLouMG+3Be
X+mvx3vffS8+4o5BkEpvJYHuK5bz2v7diwbBSTBSD4+JEeH4PLiB4dUGGXMfxcXefKAgC5lhX6Ko
EorRUf2c6KS7nX+aU9l6BOQt3JQnC6BXCHHULSZGlAh7WYouDebIxJATmLDw+CpedGphBRpFy0j/
qs5rZLFsTY7GL/BS9s3oBCTozZ+fvU4uuGAJBUAIkZgZ7ysaoY4m2nka/uqvnUBAb2nx4r1u7gRC
I+o5D+/T0HBSZ71lzvB4LlYfrDflLBCQOzsl9nfxOAJnhwHg+LsuTD8ytoYJsFHD7Vdt0g1neMQz
/X430p6NGxNY3vb2/EKWAJbAspD9eHf0NBQP7FGUR4A0dHa+26psJE8ZNio5slr0vTN7wPSeMMmT
MoDb9xJnSB3gr00nq240YJkkxjzkUGet0fbFfDy+8IRA1z0WLapMuwzIZ8IlQdvFdc+flwHWxg0o
yuIMK8J7bOlmtj4Kdl4HOFFqJc/8ZXmaEbbOJQ6ZFVF+knWwy7wJOSRl+/LGWMUNh2HifbtJ3Tds
/9sArVerRhLNmDV3bOdETmh85KOA7KkEAuhs/r/JvYhtqpxPyPTrlEsFfL4U+mrX9K9QXLJS3u3M
rY7kEE670vlMEX8JoA9Is6sZ68w66EJWlohB20jz95PfoLAnWT4cajJXGEGp+viuj55Q0ebwhS8X
E3QrxBzIaAV2RgCkI3kvUbDkpw+fLt6h/s4R6FS9heqX+fPY8I7ln3FIxl/yOWU/H6b/5bHThUhD
gi6pETNqceOXy4aIotvn+CTWfWm+lCF2rMQwrP8GopZLNfze2Ma5OzTKfa7roEAOr7D+K3XGfBoo
wodWJv81toJPA3DxpsoHR8jbF41EpdsgJuuekRERrZD8RwkYhxL34W36+Zsg1RszPK13Y7Kj/mGE
spobDt2g7o/6eyPOH83bRKLic8R9XWpJk25/XtyQCMEq1+3c32MRvXWUttiCifVnMVdrWuL2tjpe
jMoSTO0FaalpqXF9hiFWOdy6Sjwmx1ZdgUEXbCWOiQ1KRC6n6e9rPD8fMchvG8R4m81A6d9pG8MK
IplPdNAZneqXREWpMn2PuefkWSXfBV8csLN3N9uFTd+Q2VdqP6RrLm4ipEfx4jrydY7yqYbNLwmR
kXSwAUDG+y8LU5RY+8P0jLYzNXYmrYhQWy9kbUMAKYw8Buf+Yhw+vkRTxXbH/ByxXMgzbN/81FNb
Au84/oVYfPFC5phsP/wT5g3fqyjaW6JFwXX1lZJGKcym1c82nt7vmo5AtjArW04ekjmZ4T0U7v5U
Qr4yCL+OhV+5WpiZ73fes+B0J+MZ+VVM9D9nbjGoBwRyBlbFI9c79vq6FFeyoBf4UXD53Dq7/+vy
UU8rAzONdFlbtTeS5FcObeAU7nWhXa56dV3JUfUBIbzIkGG/2dnH7xggeTy34syciZto67Sv1cJu
D2kU5zwzMiePtHSJQC5wTBc17F8Qc/nXwNcL6mKeWMoSGAl/OY9BbgrHpqGYdLko44nilART5khF
OjSun+Ucj1U0BbmY0xL/gwpi5R9t++MltldEthtCH9i+/fUfQRuwMKs2tA6BlrhI+KyuI1/RtIVd
EUQTwUvLfv2ZuJsOkrWG6XE9fL/rjpaeXvV9At4qdVvAWUCpu1IDpHWkBqWICHx1hfVVTJIE2lUN
DG7IdE3NYv9UEj8QjV+MMMuUGkNl9vKOYkQAYgf/4Fof9KSjhQnd3kHYwP55+WfPCjYoZ6FdsFOt
EyoLcpB09VjOuCnCLbhAZVwuAv2lfqI0jzFLhcpC4Pddwdg4ykswnhwV/V6zwLyxFe1n535Hrfff
97PSs1C045Uj32mm6dxYkNUABX6LoPxEW9K1ZM9cZU9eT8cmAIXSNFsOtn9Xti2rHQgDDn7IV/MV
FUOVqRUTEv/DqQRkYfGukcTbPGoFApjCXKVPDUj9kkJ5tEi9uedndDx78fqPZKIuPbHiIAE0SOMw
2XlFZn8A49O71d1QOAU1Wi+jB6y191+DLN688/qEZKdPOljq2rFt6VGgF/562J5nWfmeB+LNvT6m
DIaarDiGMEkwbXfait6Ke0EK0PEHRvORIBFaareOgp8pulL6miNWXBlMudgoNoHD4l1VHQoKQY9m
h66DquqeukKi7GG+PCOk0U0/qZK0NK/um9NJ5YjaOv6USm2CN2jv+1e8yHIspxxEiDzlfc2bhiRR
/WYUO8G3LZuBf+nddJGYeU8SeJ62AaxpIcaqxxXEcqfoa3vHJcP5rKSgETmvo3SxjtEpHnMGwTOS
EsGZldPZoQLZLLeEwbYG2TnTh/hBDOPs9m4CSAxz07MGIs99KoYfOyjVy95kaGZE0D/7XXCjaAW+
ZOEHi2hk1a2/9WXXdNjDhBZ3aIWJBh2wFSQfdItmpGkRHXIbEvXkGexcqv34jnFygUNHw0SQRrg3
NAq8c1/c7b4ymvJGQFBCreMY/+YCrGZ22hO784dSnHzOajKToqDijGXP1Y7FpVVsNADWBDuXcl2z
3kkAWTniCOUbOhcDwuYmZ+1nTY5B2hr0f6C9xpCO9HZBVLP9Y4pPXgzTEruD8IgnjFAiJEft1LM2
rnqNb9y8A9Y06J27rDMB5uo48SrdXg6lwjAjWi1LghVqt0vX7LGIJLGN7+sxp2TuNGw1K0owMs15
Y+xmZTMl/JIiyroCM/9SHX8uHobcas+INB9CXmQuzKxmJ66jSYocn5vReqHf/GvcHbtntA678DH4
/w3CqX+vHzHm89n07hC70n2kRCiIS/aWvVts7cAYjXTm/F2ViWySYFwhl5qMZQT5lulE3rdb1Epx
+Kr4v4yAQu/fj3Mgba/Bznj90zzkMeVy+xJ6rwhuxPmIQQwHPNIpd0kEw7+iSI2XIz0gbLdpzrQK
jJah1Ga4qhs+zgxydTVKjnBfnlawYMOb/BVpcdCUjxExVFZZDncVqftVxzsjYOWq9vpf/N4wsA3c
oYOE8Dqm6R4WxuFX1y3TVZ/CIgPkacifAw31JrV2etTUTqaTzKPKw2Tkgd0rUWFkFz35+94ecgCa
uoxvvN7yLNxRb5+abkJpDofWTfj1mJPuptpTYoTvaFiDC96DxiJVpeLLeaAQROKe3IcbciGr0Nhn
mu/mmCWFUnS4D2HvYsu/k/U+HyKI6sqauWPrQbRGjanXo2sAK4XXAI9FFJqLpwfYM7EPaiear546
waJed/AT/Xhy6fKMVLtc+eEpL1q9KelrYUKAa2SImamrnHJ3TLq5Ja0rJWsjELOCUfWKPTwYN/LZ
Wc1EGZ2aTPZO+sY+7QjI85r0+juQRKFeMTt4wfegNUBvsvaYLus3M/A68OWKTXKNU/HiKNnQ3AK2
vw4zsQQm+QqtLNQmjbCwSXN84zhziGJzTXO27N2jr9SNQrI9BQZBvTT7xqQgnoEmEVS4j/PnsdQT
rf30SBgvXfsW0lfod/UPIp+DPJbqajylQdTdhSsqdSLCWM/7VEPqEsub3g8Yxhj2gwToFmKhLODy
a0KhIWn+dOFsS4OyM2FenAfXMgHvHUyV7mXkkQARMvhaVHuP2qt1GquhHmQ2dcpts+a/t57sPkx5
Xpz9UI6BMCUHn5I2we9K1gKxfLJwfauyTBOrA4Ne5HxKkw1H5KfVDQkKL4hvTdf/lGdz4s64IPJI
BVQUJpkL1t8qgShNHzMXcGtsKlAWLyYTua0jWsG9qzxbwZnZJPPIB9kPi197gjN6vPvsJNr2kJyd
ExDHnMgThHWcTDytpIXtydSSe6uJs6yti8Zug6IeK0Z1wr4pKL8RX7Oaqc9VRKP1Tpek/JEQnrgr
VatpgR+c2oSSR6BPnPDuEWJxQzryZg+iJ6KLJlwORuxLiJGWxjNWMvV909nzE5IidT2+j9pGxCXm
5pLmaR35z1xkfWvVekV8D0tDuXQQWzIXE75OC4U1OhLoCKTbWclpv1wHS5zvJyjAF+3zH1OMy5xc
1osHpdpWIdvulr2CeJSZiuw3VDRzsmXw9+DxlUra0uaH0rigGrJaKi83lclLF5Cp9/Pc4X+He+dH
bD7eL5Ryryfx7UbVZDtZL+uu06iRt8V0Cx+eaRUv+fOHp6irDMGsxHXu6zCofP735z0phrjGImlX
qpmwlkPPo7mo2+j8WP/xW6fWz8XQN00D/ynu0p4J+wIUCKXOQLarSBcwh4emA8md3Gnb+lC3fhr+
4nGnQy5m81r7R6Wy0Z4NsWwPEQUD0EoMTkMpLQ8G2r36BUC4qgQN0NlTREmKysCFniPcvk18wdKZ
x1pijD7s3QYs38rvKm8WBaKoFFc8/O8YwhKdP/lLe/y8arwUVk/2Kiz3Vj1lZy0Qu2p47TgP6/6H
rS3+1Qwz2fqwsvs/cvDQp39gyn+EAG07CwyfD+1JNrwghvi0RdMq2PixqXUNKqJ1LTme1Znae/nu
VLyOaIcWmpqhCIDPamoiZEExaGlF4TZtGaX9mkqFpk505eAVUce25QL/9gBi2htRgF3de/e14XsT
Eltr2lkZgrZz0JMO2uxx/vSq59SHe/Am+DmWe1XNmrBwFbMxVhWhJhSqLTGiQLnLfJafztMBxkNv
HDMWNZGT0wxZCbkRWtN4UmhAwZPx9eXC9xQnU2f6kFsNJ+/oFMZCdC6f17rbmVLCsEG/uXTmZ6qS
hsfnPXIiyI4Cj7CwJP+4pzxsj7Vilu4QGGjsHsT0W3ourd/zlvla+9kg9Mmcxd/AycHGx+mQHYFq
aEF614aFad0+3SeNRfdFiupq5JmpR3RvLzu4xLYcmvtksKVhlTOpvWniWtBNe5t6N0ARmjkHZ+uM
2awMVNwsTJP38QV8lEf8CGpdO6w1cYQqGUZCSC/JEKvB7hqc8r8Pv7QkeJBrQ7a8JtQd7BV4R30M
pHLu+JcmZX3bmPzgLHkTVdK2ntm5hFSmnlXMcZQPVzs75hBJt7PFN53zu2XU2sBeNqYqJyAYUyCx
RtZaHZnfd8OSO6nAxb+0yQVQRzRrYa0qOZRlX94agM+gMkd/KezU3KvdQ14n+D5EqLkUpt5stMo9
+J9tw9Ayr2eUUylzzMPRG63UB1i+l/or1iGU8+7Ez7UicN0S3acA1EDSudR9LKZj72m3FrrPbXMo
KaXGYtBW8p0XgMmOvBtwAMNWBVfcRkIgjBbb11U7hRihvca7TWA0PFAv293dzwf+VUFhoRsKCUV8
qP+qFYm4TxSMzqZUPMdM3JJFQs1iFveddf6yCPK/VKum6sIiTXWRXdYFkta1sW/QiyWIQT2QbhtQ
rORJulfYsW3/e0bfQW04HnL6Z7WeAAtFsXFuItyq1NxXYHLkoI4P2NLYpSuhH4svEKthQbIdMUug
Lsf2ckeGz3pB+Zif5LQaO8rxiBM5batJdcN63bwbjNTK9xrWdG9K6cJxAuhU4Elo5gT50kpICHUY
bIu+PtPlMonPU2zD2csyCqYn4LrFDUvjKIjTxme+jfImYwpYq1eTeknxwXmtuBqanY5D9Dfyy/bH
433Ctl1quH3gpBxCx+vGSUvOFh8Qk7sFxKJ5Ol7ikIgmg3BNIET2Z3Zc5OJjPSdCoxksfPCGqR7V
8iAb/1Z8bqY3HCDHigFnFHToJvwkOEK64K19etOMGp+JNfz2WYIJx6gfiT7Ix04Q2XeYcb2v7PCg
FMkuYJa9/3jeGGltCDF/6PSYQ762UFnLfHRJIpB9d/mRPPfJulXuWMZa3A9vKuwTm1jISvqM9rwz
O30ebo/uSGNWTgFNfcpN4OxYIRcytOy9tLFhDdaOMoagwpKttgSV7ThhmkOiE3jnKjR5zb5UTv+3
ZUJgeXSyPRPuvjWCfOZokJKhs4QZSc6jiBeYE3SlG3ZG/aGEnZCegYSN0gAfPxFgeFyY3CwSmA8C
g4gtllKoDxFkzRAutPpa/0Zi1flLIshhY+KVr/gqohD2/QwBtdlobu2mSDhsRC1KsKjrJ4nCYHTF
gVKBDdcA5FInqYGYGGH/aCQQZs4Kw06vwygeZRNihYru8jLnGOmPmGoNf8A3Dnkk9UqhYaX9LbVo
xPLP/hb03mvoTBlkiyiiF0B2xm1AMuWFD1A/4zw2eXZAffR0oI/JRd91U/aU5hKV7sPnZFjlDq14
dva1gKV28fPceB9spXocPHPnFfAMPjCHZ4Y+xy5rraR7935peoSQImYEyH94k/zx63Rd/PmmvCMo
Gyr/TvwTP1TtNI4Y+WZWRjB91YOLsdaZEvDrfCRIqX8YaVyrKtPvQgA/TM5vvZWMPOd6NsErxnRY
/PFA8t7FfxCZoJgkWG/GHQt4OiP4xIBVHkJBm+NJmw584bOAWFmyxS0ZwOGQVHdT8Zd6hsRa+Ioe
xcsZnsySQvF8UWrxHyfiVy98io1X4NCH17vGe9RqNWMABgS6KOO19fAk1eqMVoRRhDeMQT0m6y0r
L5mNt7eJqMe7rxvlAQuQuUu6EC7N+ZJsd4dxoN1DgJVKE57mgrLsWmIB474Anr2bZe1An21qP351
L8sE7wlqwmWUeQWmOsoIOLyDOtF908h3sONfEsT5ECfwAEzyDReexTdPuPmhHFyKcjKtUitK7Sv8
kwgwJAIKkq1gDtrnKjALBk6pIEoFvTJ8tQHJ4+gINRoP8KEV7KaiZRng3AcFbNRaI2d1Lwl5f510
w45sheVwlaTMmY0LhPIBH8Q6QINl0r1h+voHs1P+SwTSgLlmbFqguNkIViGZu7apcYMDakX3j0H9
PdOhFXWDf6mw/MVwZiYeLUA2l3FiQOEA7I8/5OmN89wNh1h7JyeHuBixS7EFrly64AZfjsP4QGYQ
tYb5i78+p49aNGX2rGJI1VdFPdG4FatTJDDL+hllgHTs2zX5cRq3u9dScBR19sKqMYWlPh5oVszO
UCBpphXHlvlntNmQW0cAisdXhf6CG1zGerOUkX2HTxnvRBkcw6MIEBou6fJnu91x0AohYtxgai+Y
qiVHXIe8eG5f+yREhxPoP6Plsl8gZLfCTZWiqIH0sAw38H2lLnlAZQ4D2TExuYtzvtPuHto+PKrV
g2oHJR6RwZS4oGvTkG0DpQrqkc1jCMt0CmBo/EaWcMiAh6jZtIvYxgjP7fP7CA+x2inydglNIihD
JF9iOHr+oUZxyngaybM2kct5UnSNJMGQMJpIZDUWMJHv6PbFJHeoZ/AsVVd2Dvy/y7iGgs/HQh0+
33UJjpAarPN7532PaTOwPmA3cWT2v7qzsUMUtiQi9dwbPPk0PFS41kXcLfM9WC7qWZDZA4S80rya
x7Mrjekna1DKIs/viHtHEoz3QhQCMQfv/akgvlGNVxsOYbxHl+2MnsQ+xqaZNPSNnVdg4i365Ukz
5z2R/FV0pOdSm9mWGMF82mNWGM5HUmInbT97+APQcMNWKTv2eFX4VEYjTtyJ4WqHiBzd7ZEbb0Uq
prtwHJkO+3J1MGICUwxvzA8hMLNz3pIeTZNqqNYK+QjBGdw0Liuex1ETXs8VNeWAQOs2lrovt8jQ
EC4pv7xrEph72lGvA4bXifVxrNG0sgXTQuFh5CW+A5PpDxQzNopELskm0b1c0lmP8pVzj3ObfQmy
q/9YKAHpy806jlOjcoseBqi8nYkwJK0NVss5W3y88aBRmeY1+9nevoEWlm7zQAK11ntz8lzaUnK2
pEduFTnC3lkEG6+cE9bir8X2P18/rOrvIV0HNV1jZW3O5MKDept7wi9tTeZEmqDP6rH4By+qumFu
ycjDMJf3Pb/a/KILxIC97cLMTWmE8b6elxX0oIWtOsB9tzxci5LROIiWQxn2WoDzwDteLj/RZYVu
3lBpin67/hFNYZGx8XJZPdZJdu9pDnZcnqhzAzp/JyNcvVn33gpNdV4wXPIKpT/D2DpkYmpXDjbt
g8AFW2zsOi7Z+Lh/QOYiucj/f7nkd7LrZYw1HnSPfMqjXq7ewONm+U4/1PNW35t/z9v2rEsf4kgy
hOsOKHf6G6y/F/4SIVj8jKCyXEW5Oa9ogUKoiQzHkkRkBHnJLXD5hYtCCLIUqB8D7rVbai4zjQ2S
+uNQxv2pA5kOJzMJh3E93unsNA+F+J7nzW5kLX/TNeMd7EjEccdsMm25xjTaH0cKtjkhh88jzJgr
xHQLduV1i35vCU4xmDAShUjExJWYdlsRwmwrC6UrsIRCmDPWOdOWO/O/N1xeN15PJK7Z1KLg4Pgi
rR0+SPEQxhSk0nnsYBkPYUQxtaXYhyqb/t4OAxERjC33GEzF+v/UkEyQcq8gAZvsbt4wzvpDfU+C
sNHtk+EGKnoh1HlbaFyNyFx9sdzfWjClpQ8n/lQFmnOmH7fZI4d2EyiBd3+F3sWOT1NAKKruCLUY
wtIegLO/Z7xLRNdczNmJIyAUdm+nFAwmSvoTM4bzcjQIFQVkZmVILJUb4BOofapJHEaE5C7oHf8X
1M/ygwdH5QivQwuy2ARQ1zgljeFZNsb2lxTMqPwl3fMdyfmCoTKyWsTDBudpGGbZ+SQ0oUfdwgrf
AVVgcnIgz/jiC/cfQ5bX4UVIUAKy0s+lv8svK1S77V1fMg3k39VZjCqxW62GhOqjF0h3Sk040iB8
DzOOntAslF0KdSFspuvS/vvRm5H6EUXO0DRxmTeB9o4/gShizf4GMwbDnyNZKIhgT9GyNGs2oBbn
5t/gh6mTbzD5dhbbNzMeNfh1Qgi3RjteBMCk1UWNJeBuk6Gj6iXOS1FfhVWqJuJQ9cB/DXThQIHc
Q4Q7Eh73Be8lgAPnowTAFt2C3t8sACvWlL6x7uMoHS40Ntin74RSkc1DCYcmHh7WQO7XxZm8YjkV
6oqtm0gaLVBL5n4PeIpEwBSDEgMKrO15DDeYsuP0sUlz20v6qcK0f/Bj2vwisOtsq/PtrVYNVzlr
FzrpMP53sYPiIO/Q8+L1IjM2+smjw+0V+KwAP4JlBcsPnmH7nL3HTt/17WbcvDVSIHniXpQU/8J+
+yIXZiN6lmEZde4mGM/PtLCqPyJWVOIeLQCd4qNBTx36cOJ8WqlfjWDXIFBUDLNTIu+1XzaN5HBj
c6m6Ppc8D8oajYUWldndBULSGA/IEMUcC3oAZNq/RCdAJaKgxlj6NWAWx6rZAB1I++iLiyaSQ77W
fdUI348i2/xi0RGiROwQd9+wzKSmvh8gaeir1Ivd7NIr1luSEnAbuYoRjh150YqeX4DFKSXgWGvV
tFXvuA61mY9CFSQimbi2KIvCa5bzbr1Debow+E4VVSYPLTh1qwr+gVVIOkqv813u3xYZp5NGA8Nv
B+uG9YRgadfbxse4x7i+AvRWwzzA4RCKwIu6GCmGoM+Ox9M0gsVvXfiCM1uBpDpE3rYqsjJxStm1
kGNrwkKK5KeF+rF2cArKtPJpL53V+Fyxuqs4yLgRCgBexK/hBgSQRMeXO5vawzmCzLT0oNgbNTNJ
a1zeIEY6veA/Vf9+pO7zarLxEmdxwIe0c7TdRNbZVele7oJ+ZC2mboHlL3dse/afL+9M1hGjnJg2
ZX/TFt943mLuTPh8ZUyGyrep9Z3f8Oh5+Z/mDL8aOO0EjtWiE6c1l8RR3GMXzpNUY1Aie5ailyVX
Jfc63vLCW4B7xXRdNLVRVncUBpuc5DTn1KViSK3PBG8NGiPP+PNA7ivoaXZXOyBZEXcLb6tIXe2n
VACPDHG13PtYkWcivoCJPkDIoe82fAwqR/HZJUaLuc+OK5sXvt8PSaBF79bvsJwAkjtk0t2gpUc6
ifbaZf3xaU54cGxDosyMOQ74wR0T2IEWZrJRljjDIDzs4AxxcmSZNEt0a/bT/awYkHdgQsdFTBRK
A9Aai/TtJWSIQBLE0JIxqHBNkENH5gDsfNJtdx/oAqn1nklAPK9mxpKh8YH89mYP7SvhlrX9ntMt
SwPmpZqD6WtjYmSalNiOnFLh2RKN1Eh+crrCvLcBk6ei+YU4YhVft7YyGovLLHuAO38dM5O/6yKc
eYPl2XHBZFFRPQSlOvyVTF0sRQ8OVIavvBDe1S8GH/nPW23R0n8jdkgDrJlN+UIPmPDZ6o+NfT8A
4ewiLMDTiEGbEJvtgpW+1RQtfh1uQOsOJnBF4LneWyq2MGuGSmUIuSD+Z/YG3Q1zYyaRet7llWbP
E8z9CI0BeiZQcu23csPFr409jZUHhMc+RtGncY5dC9tH+0QGF1Z7OIo4dgLorseqfiPWRjXKYGRZ
iPRjMbtht3wkusz/YZxXvYp1nAtFUzIWa2gQvBAMf0xW/zc893FxVGn5E3Yq9fgYU9VuYSkjQ1TH
mLL2y6MD8v39mclT3O1pT1guCU3CxJgn+4nDeI76d5dH/Vh7s90YSjMpUF4JmnW6yH8RgVV1DSeJ
xfHM9YbgpEvtX9gWaCNvdYxAleoch04AS2YMvDoI7Dd4M3QQQaWQbAxTKkNNXk4iyg+gvCeIGT1P
NT9hBbNIVsi/zK/jeqTKN2hQwy/Ni7FiIYxP+I4FsA598G7Pmed4pFZY44lt8KYoX4D85LrCuljD
KACoN5ssqnFnNoNRSa0ysML0re3bzatuWRyl1K9w7ufw+P6yPAqyl2v/i1fVZpjopybe/Ee4F5i3
PenaPnaDm5tKeY4WPQ+mp3bY1eDzlCPtnl/ZpzOIFoPPuSNMGJ+QB0UoNKnHAlAGT9byxwqnjmb5
4Mz6QQPTipCBuI2q53DzKUBtswFiBT6dSASvwKC3TgrJby0JBQteJkPppvQ1qAWEdJVDy1Xh7HYM
hsmNcvHKFYFpIZeONqU+lkdGIN1dA3hwMh2ljIE5vE4Ft14ct9i4nSnhIGb+xlmYzVdrFXEHk8Gn
wC+piBL2xhHVtPg9IY1nKX5LXMoYObyqBUk6EUGtWM+jgDkhkMatcmLmlao+a7V9KJkIcUwTplIy
rJSlRghzOgUqPXtLE9+v5raiin2qeAoo0JUeLJ0uNnwa/Dl/sX80uazDDdJgSWkrrADYbWZ3cBAz
LZfwDrrdOi6vHfS7co/An5w8EjJLoafUf4PBRd6LhOK6eQljNLN3ahA7o71SnokhqMFXGAfDir1F
mvwWyIwNCzlFE03OhtZXnoVNExxpNFznwqOnsc18Km3mBi955/NqfGIfVmxMJNsk47waXnwW+ZVn
MbL23LOAzgj6juCzjVc6fQ12wpXjaDtUunApDtN5S0yvqP0aLlPttyUv6YP+zszqrkIg6RHyIsIX
7kVda5csyLnr8Er77uVKCCf0L73QP5lrlkrhhRaDnIJUg4NOcdMbao0jLU+oP9y6LtDpqhjzlkcd
UuoQC2QH5o8M+eDHKQ3EAtkp+ci3lD6CVyZFJaW+kCDGHnjHS1haRbJZon3WRhR1unXcyHiq0EVJ
mU+Xbyj+ZYTgMahqXlGd1xQu0UQ6dobdzYH6HMIkwqcvQ9hNBONDnUvqMkVz0wTci5Yp+AC2idx1
Ea5Xbe6IOMSRSrFnyI5xM6evzCNmEYJETnLgc4iidUEky8WMHIZXpUrcUIujVkfoGm8leAeRnCvr
xqCk57Fyqtm/gWaH14hJ15GdCwSV7yPHZZCCvJVqVCPTo0IDFuq9EPmUi05pWaIjwA7PSNMQxyzv
q/BaKMRkM/uaRyc8O+1naNlS51PdDVVmuFTHLWpJqcuw8e76/NLEXczTJgmi51gW9XhHpnQdiRfI
rKlxVElF1/FoX5ORAWEZeEaBTJ1IqcU5H6LN811St6YVXo1IpOm+M1t9/zEUe+rFqGc3+VjnxymT
zTvZKOKssw4rkSB8cVu6xCa2QcSX3JRbfOc232uI6go1vikR8mU+MYkz1WnBg+vGKryapqRCzxXE
qTZBuJhGuNFejeqTRJXCvBWQ6fo8BmFTkk0+pl4vXEOvpLh9Z6R+kkIQ9+5aE473f3eh7CnYIQun
jaEN77zOJNb926W+Wn7GtcR3FKj/hgYcPukZf6TzRoy1gQpb5vSrtPttlOIR7oNO2zIFAELEVi7X
j/Z3Ewiap897Wq2ecMC1C3WvMfqZdTJC6zRP+LPw4thElAlqLDMPMKA06SEwBzC+Sr+GBKxYpHAQ
sCdo2DGCthB4JHPXOMD7/PnZUDwu8caOzIOKb5klCcDOAY11UpTVBtGxDuxTmXHvcdaffsdVjIct
VPqQjOTrHT86lsXsRJEc4nYC3uoRVh7mSNPNL/4ye1BqCWkA1ZRtYv7MhczqarLncN7Kc4fDxL4C
pUaa3g5rK+XH4eAw/nzZ6ut/+kpSqd1yiyahuBPcJ895V0ZdFI57uuqZz3hvTjfiGigP7OJkL80y
5RGTylAyRhq5zw4h7/m1PxDAUh18f+fYEuLJNOp+82hJ1kOJynpvX8dWz7xi57QqZ1qjyUI3Juwp
QjW0UV4RBqGEUQa7Z9g/8JleuFGQyiB9wJanYH1x47bU/45V1N4XuroOvkuekDFuFAl3i9t2Jlwd
Mc7/OcX+HochDP+JRkOCoWPx7+DUULWTxgxjqSCZPMhGlajnlcHbPmPKocidkzRXchm89XSO3Hxr
p81BTGKh9latuoRu+5HNO/2mVRh8p7d3aFp63SVnEERd7H+2PLyBenw0k2+0IgY6z0Lxt6rCrTuu
jNhpJOHo8yTmILiyisM8e3p6n/9cJjM6SDm02GdIfGK7S2yS/1Mt6jCKi3pb2ghEl9DvUNcMYdXB
NBQ0VVANUa1gt7lzbjLg1fH9dPzb5EfquDEOie14mllyj/bI6Z8FvWMcyex9q7+5KDmHPMpMktpw
8GqvQucGbfzmYFO8V+6tuMhE2kLeoPlDs0PzZfLidzZJMXWTaZ3HfBqhFtFMY+9hrzhr2iaYMzci
zbBmozhC0km7CY9f5Wpewwdv5oLWkCSOgk1OuIml2DKD/FgQecqFVaCtGwZwIVofPEybavV6bVud
Mide+rrupbAgLahtZfuetcjZQvozNmMAywvLy/+ZuzE8a1HVSKPLVwOcWJC+3ljjSbsOr2rXH6I7
/TwNrcriy9crqhkVJ/Cgw85AcEzzwyH3mffAwbsKC5QHJak8Rwu5WXknCsQ5HkPD96NuRG0Pl5pl
29D/yDfH4LH4wF17p9k+S2EB0562t+rNCxgXHb9WGEBOr0SJE+of3MuYu8gFbJvXnAJcRZLd1mnK
G0L07P6CPDo+8aM4sT5xIPkKvslayuJojv2fcKM5xXbmzGQPsZTfAZKOew+ausNKT4lZNaOq5tle
8yTqrjn2DvkK3pEkV1xjgZvgUM7ZSj5r5EPi9w/o22mx+Z6JanYSnaRax2BR/WJcXWMUItftIGm8
EE+lNEm1eIW+bSLkS1ncFLIVtxG9Wx9xhYD7n1K/MqfZRt3UOZbk4rhBKGlOqgN6ujsmz3SgCoEV
frkOoSiOVq8LRe1RAXGkc4pAB/ncOkwfcfCsjtCbm6vBC5genz1mTRBJM2sDvp1QLxz8MebBTBCs
vR7+CcZOzpPwLY4l+uMt3weEvdt1+anXH/1H+nMwg4Y4JAuZhVBQI5PHEAYrToF7vBsF7TIrKXmW
DA1uSDP2c+TZxu2vymrxKUhc+qXQttvy7Uf8JOU4Ja8H2TILUfM7gapTRUYhrNZ3fUOVuvEGS3MK
SYhYQiOLO8YhUHf/R7d0YcQTsEc9t5EFu9dkjHuXVmyArQz8vHBst68r+xCV34godtQvCKpCUuOA
j5PFbDMU9T6931c2205VFS9YUfVYHJ6UsKrf8sZOAJYg1MfJv5thF7stB5feSscurmwmBAXGK7O4
AIgpGWcAExQIsEgDUDPXjgh/9MseqdRihc6Y8aiGGoto0TIsUOAg223FtXpsGxQ+pCuIaVWf3vbf
AQdTLW/5vB2iMQQPyUlgSlMWRSNfkAD+7XKgKLLrZIbGSQoziY9YnCftwAzvbYJoYOKpkku1eDF8
rifpm8swE9cBAPwy7f34mQY3EUwuaUK9YXcC2Lvh9UAs1sa2QzGf4xFFLCjEcfXwQEyOCnw2RUQb
SzJ16Xpil6jsnrTb/cX7McdgB+9MwK3k3YoVcxokwVIGdoi3nZsSOsC0j66h2OzEWD0HXsteLQ0Z
2ixcg/0K/8CYr541JUx9O6JE3UrV/ApSfFHOhxZ9sV+hh2eW+PIeWaGJxz7yvNVvg7pkDySoox+G
vDqAaYErLhLG3jpgP2LHjNxJAWHyWDJqfWjoU3U+Vl0Fx3r/b/9rQPz7XoSUx0BeNap/sR6iJYIm
jzYu+I8Rb35ZUVGSDr8w32S6NGYgzWSsv64fon6U0hhFs1rSmgxilbphiaN+/AN9dkglq6rXI4Iw
FrwPisyXxPLS92H+9CxzCzxB07+gWQjYGR/of9cEHohqeXEWx22F/bxcWCta9Tbb/ku7FpUFv9an
fR4SrjDhOf+ri5Z95EKjREHl4b9pAi/BN6Ru+dFidqihigeCHCoUJ4IvW2OtbgCGLRgOqX/KkQto
ZnKaiZNOEYM7v22tbGJe7WID478Qs377FRAeAAXUwAujrqgRt2IWdm0Oo+OxGh/FpI1QZsM9rORx
bhUIR2NLb9xhQe3Eu1A24I7j8c04Ux01kuXpj2mgKqdwuMUVgGeJaunXx5LJsInMF0B3lnolfC9H
t9GrJVNr9wboC4Y0t4OIfDuhU09YK+ESlTPqt/fZKPZDjKrvO2tCuF7Z1LQjyagOh8T2xdZaFo7G
zqLQUnIhc9reofCdSzaN4PAOfLkQciepyYSNTtXTCs/n7DKnUkzt45aSsef+ZZ0L/K2QEADEgdwV
Wg5JANptik3e3udlF4xWeL8paCZeVIryOKDdKfyTJ5F5B5/j9bmZhAYXKqd3cA0+CjHPNg6zOtET
NXAmcfC8pttYuKt50ZnzBvsQlgivE1NprUSIXOYB2MT6OM65ed90rj4EsbXM0O49Fg44XC0epwn7
BEhQ7jOhVsggM2d7Qp3alp2ft0sIV5aXWVYr4iFd6Fsm7mJY0s0wo+neTJDstncYpOt8C/mpu1Ta
GQZKG5N4+mBbDz1Lyjy2yvYKYuXEPOO749JSp/rtwVTtFycPpi6n/O86GlCSse9aMbd5nnL+8DoA
xbhtJ7NXEUQH7IHqcHFY5NYrP0HwXp8Epob2ePA8XZr23L8ox8+dnNSPUND1S+oYzj8dUUsrX4Gc
jvyZHOfYNZFmGXYL6tOFj2cT0JalBeXU9n3hxU0pTPu3AZZWd5zFgfo6bP8Sw7rRiBn02T/nS6qP
Ww7Lui24qDx6LMYOVJbZ3AYeWTRoctc6vWmzN18A35qjVPwJVzrlkEOAyHW13I3B7axGB+QZ2ncY
VEvSDSWF/fIpUDGR/qi/DDESp/uJ7nt5Egi7Ar/yxg+yKnMKGLD953VZFiK+EiQZRbnB1I8ojrKE
Rdl0U61xXOUYggxWMsHp/j/PbMkOkFAWRVA1HRJTFA55SQkJWXl351FxCZuz5JVzj+Fj9O2uotaB
E5E9Sml7My6s/VzEZmj03if2OGlGowaPClzDAnl2FW/2r1YRtSxZrpL+L0+y8a4HyafB6GPZgP8v
7JBh/iG+aX9BqBn8yu8zEkOTj403o/ANsxgCcgSWeCHvkQV/Ceg7ld+6WbyrUlKRvOiE8EzXPQPa
D7AgCASiXRfJJ9ZsIFEbthnakbdLXAaWreCkbBy2HnpVyHawzTdzwYk62LJfuxTNfQh1WIM2Ztqx
JfORh9hC+4AGsSk/qhcY5eN0WGJ9/LEOpqRpydFTbp1U2N17VK7XJSbIvCG34VoGkhAp+r7TgAKT
uHqpYRWnaa8HOBrtKfZJjVOF882PtwSefRnupfllHFsy0nR6wcswqqG/nv2jomM+vqvjvofhXTpN
bxmgkygdbKLYWlMu2hx5QMtOXNDmHdA6MxevYg1mvKrvShPKOjnorcjASObhT9gfbYs89qLYU35d
Db9Gxu8wSTnaQBdAhM+DW2tEVN9DL2MX/5Xa3U/ShkxNjK5hh0hZoC18abYzPhgAtiBS94KRZRiq
pYXngeKJn763GJz72+JVSUpgr9vIqVUn7N+EB4mdc2ya6ak+kvoH4Ul3V4EdQZbnHKHjY1cVGuRn
73iZfc7le/oEQIZrICj4OTtHM8+6ip5L3xjOLNCJj/3VQNNLjRhGTAi7Bphmp8OrZlwhbRiT2nw8
2e4qIUMt3XN6KA7JxPdYXaF9SppxCFUxBVWi9BqLQRZK9DvbMIk1DZBZPlIydsNXazTafqgzNhAJ
kFEZA5nj2AF++r6hNz6cFokFNINKuE/HhSiq70h+UxlEH9ITqyNgDhaAoEnafWZaCIr+iWTjKHbf
DI4v4Idm+eO7meut6RGdgdpFhJdwfdXo3GgH8g5TcIdZ+198pm0gtgYoFrHvNBCLg9R9BLnHgl+O
bonsnFfJ1srqyRLDFlhz2GL5OeiRse7pSwyxDV+jLSt2ygrr9qFdmQ8v7RxJsPrAVSe9/idhrlRA
96qSlfAOcIaLCSxEGWGnZNRDf7obPjT29ZK4siR+dLfb08m5xnyqsnJUGfmV3Fk5WIg0UB2cr+dV
9D3RKFxMVbtpaJ61nuJT30azlIiW7+sKeccG1lNpDmtKtYMb+lwGJ70RDyd5gT3dF3U7LUQESEhZ
XIxl99UP3kfFGLbW4zc4Knm8LrdxKZ1ZUDmaysgQKqezVsb/1Anwktpko7mq3hxYJEIfrKd+MeNL
5G0rtFS1RenNPl4DwXKcQsNL7xpaJVMGHJGCuBxwdeU1aOjWVw5Kd6sOHj5tsvmNgxQ3y+FcSNxi
ApBWGJOSBHcYCXPFBfq02eg4WzbPBud6tteus8IC1qXRM4aTNcY8bmKSMWI7a58t1eomZQLqb3tx
LhwweQBTPXLx100wZrmeItm/9gMthlfdkIu+gxnWypcwZxe6gJ0X4DfcbqYOOME1UkNps6xIJyhI
L1o7jEyL3y9brx0acXGK9JHwOS3g7zhV8wFxaASa9/H+cIi7vIwEutH5CQr6+ovfx73+ng8AbQub
F7fyP6Fy41ntrgpH3SJjHS51mcl03t7On0fwOWUbZMxffsq7s1WLhixd3KvA7SnXAygVkNNepFVM
boADitu5CXClQd59fxoh1jdQ1CgOpIROHBnKtH4nlvL8gNjMrTF2QezN0rUm+EEM5ZQk+ZIQjqu6
LR5SA5/YoT4U/pUDXYK6fNcrOJ2JDD2GWybITVh34gPt6TI47BFXraObMh4DOZyx6uFRMKBedJdQ
T8/G9rmPdP+FlUTLTyGFEuCJJM6XPdaAIyJw/qd3IDc8Mft3/Q6Avs2CqhNmrYsLMYPzyJuSrN48
QsbSwRhHO/hZHxk7YlDud7TOAzOFeSwGo1wKZ/xRpsLwlKXxgo02ZhQgwTOIy2wY0aC7S8qy14Sw
qToAK0PhMsB8nsXMAP/xF+JM13F4oziCXeSpnHhtslv2yQs171LINCrdi2YoZv1IqSuY1wHLha7K
nnF698f+ZSXkxzFqA8/Abgn0pT+c8Ub3CB5XXUNjhUeRPICU0BdD3Cr062Jw9Y4LAjCsSdjz9P1b
OLlNtAjBqVePnysCgG0kECvsDCK2Ig49U9tptKdf3kUNKnJws/3VZQF78Yjm5iqoyQCVF275k3iq
qanPuypB9XJnIdNkeOld6dRRIOLsEU0kpCHoHC62bow7U3zLjviSLC5ieCwoxn6BcqneADm9gMu6
afCeduAVqmlBAf8Ez5fbXXMHrYYG169il2gWSwJ7Ef/I0Vv/L/1gBOWk/ZYwjRLK/T0Ywskoe8T0
yf65aEF4W+AbSPnByk0RGWfXkbBqWXOH8bcnJFLn87LMpaL80cftHHQwQs8KxiMJWPWiyG07PGb+
6RW+9AeYQwb/AT3b5avsOWbnyOAboHnx74ZFLwVltKgmGDXmtbBNhZDQPhGKL1Cr975ko1Tfe6SE
02/l2ofBhYYff8GL7ITb1qvevpcmo4+SkyVPz88szgtY8O+AT14gG28n5myeTwFJW9gSgOlUzM+d
5IhEJ8xx6DTzrV4QIICS2xEQSKmlnuPGvMMYeCF8C4OuY9m8xohU0Z65U1l2t+ucD4aXBS6OwhY+
RydMXVuTChD1SdgULrb5kgDZEJnV3723swF7fEloIjVKEUubcsbRf4SeGQr6j9UJgPHoyVGVz2DV
Xu1WY4s3eZDLfmljVgsSOMuoGkpowqXHNtvj2FhWde1aq/LC67JcZpFbjX7SHlAY826NsNApfjp8
2rs8BcvmPDAHpf/sBUYupxB5mH0YPsHtnBKy6M5pRryBh8+JsCZyuyxwK/pbf5Y5ngn476+04A6Z
oT29H42vZcQXN+r5/2l7Oftal49DQ7UFuXCSUFKjrc7d8i1QKlLkWgC552Ae5vO9NvfeVpcUr73O
T8Q46hOET9oLbgIedN9tWGXb/ZQcozp1jdAkTCQI6nL7HRh65HJrDXuN2i8vnO+Vjhmdql1rk4sY
z+vIdWFuUJSyegHGw9VjxyuvKNU4f7zlPLoTx83D/dOehO+2URoRe2WC3jV8h4G3uEW/3QKrU8zu
fTJyRVtinvMqmL0kk6TbjP2gScCy+Nf9RqMVLW3uXRi3fbhbfo/8B2Ws5rIyQ5HQoZYLexS/5hh2
hnTgPY2ZPeSCr4AxsQV9owSYqBZXyqJJBobIaHX/LgNpZJ9kgiKQQ1Y3jjtmtYeEbXROM6K3KWfD
juMzD/RseM+Vho6S6G+n9HKCJDl7+frxfmpcGKsd0p+pV9mj+WQ1jPWp7iMNOsFsb02o6vrOVSNn
BYQd2x18j/vdjzDHBrhyGFTyyabojTO8BFaBys/v0QTZafCvlZVkrBM5sXEiKrm7XUgqHHLjH/aq
Hptwb9/35dFZxpxNmaBfZTMmIDjOpuIbu7r3ndWIJkn5Y4ZfdTXdqW2DC8Ic+tN5VcFE5YR3/mJy
avEousbVkPQkUdBZEJsoVAQjhVRPaFnLuVuXqB+szPDlNg/u9p29eCDKGYQIMTcvIB+EnJHrmu79
5HVpaLo8hoX2NhIKi0Zev2LLI8GmMDQ0ZeQTqofKSLKjvgZNaid0IWFQJeeVJ3Sckw76k1NkMfzs
ax+WErQq/R0fSwNI4BZVsi/3WNrxenwVInMuWXO5rNbTy/MOY9+Fxk+dxa3m1jT9LsPEo1ONO28X
ZaZzvdI+pmDUJWDzHkWq389cU28ScnzIZZzP4ckVcL0UwmVXQkKh8fa+hSMTOZygENdSOM8gms20
iE0ULSX7s80EDMsHeuuwelQVm0IuGB7kVMV5Nef6MFFXaKGY0ki8ZGsoGPmz0mPpqUxPLUCb4Fm0
CN6bIWEDSrM3nJM8zMe1S+1txPPtaA1ab6Lu9Y64LWJQ/Hc69cZF4BGMWDJghCXSnTfFz+qjl94C
G6L7KQtPUEleyrK0YpssU5NT1OFMw/plMVpYACpb0KXvHmitTA1zGHxUKiBzt3QNAR2yQ5y5+U17
vyFrCrnVS1zwKjZVeXGvPmGm2x/OgjJiOljFD9YnY0qyzGqgOl8lnLmtNphPzaEdViI52SVsQ+fH
Xo3Zea/ZM1agYc/XX5JLg7dbDCDT/kdqeCgnWPYfNtIM7rRNwwWVFAbIyN6l5EzMEBlocQi0FDYZ
uI7Zv5DDGY7ay8gFAFZ7OfVB0fB5MCbCZ11BqRyCcZ83ZxRGfN1Hzktl1c9xmz9IgmcuWXM8Vl7Z
CzwdeVlrBKv2gR1BMau3Nv3OoYlr8FK+ZPvuyu/ydSvME7xuSmdPPJKC6IJG5lh4OQUtMqBljSeg
5bHeciXRavHF7dg0FG8Vp3uWphUwMOVRy+qnMEY9yh5wIPqLQYQFS2SwX4At+JytQLv+2UZXSQ6p
/OGWm3itsVhFrPjeNrBXf7Wbt57X1GJ5qOBapUIDhsSM4bydd/FVSLahWNNMRrJ4YbRSt4CleHQ/
n6oksN7PY6Bbxby6geellq3TUFCL5F9eHgo+4QjsqcxXJGuJAoKV1tr+aK+2oEDQIJuTnxXXDJw+
mo8KyAMK/B6QxyP91n88WjdRlzHMN7jcxrJjoBq+Hv1mzmKGVlOMMMnB5l0khLiSICm8fCJVhoWm
TizzW1kUhGgLM0zMSGbYm0WsJtPW7/ntc5bFv/Ua4wlmFdC5H5yrzLWbFybxbPZ3QO3UOq3XRL2f
uKVC5HEIqTZmF/RFG/ACtWYYvNaSPTaAjDXMSkdHWnscbfKx9BLQQZPYWcmwXbmqBt9B5OjWK21A
5arF27lJf5kHJ4s3lHGn+mZDE5fx4HbM3fh3AfRkoi3Q+t0x/vVBmHU+oNk+xi2qSipxKfeFurW6
NDUDOEwLvTqOfjbAH1gj3J8jBV6yfhnTHbB3EIcxhx2KYdFfclr683MMo0BK5y9a658kif6pTjHr
T+hN5UCd62eH55GT3ypmNKnyNkgOWgPfyMvX9YshY3+L0e91c5EinydEsWmPuNtoFmwrPBHbiV0G
97iE1E0PzKn5WvVawFsCUQhSrlmydprgN4yncEexE7ky6mmcCuw0Nc2ANoi8RgfXv2Kb+QtzjCnY
fvn+pagnY9fE+r0BAKb1AQ/XhO/IvsOdxWH4HtPgAfPf7XYyJoWHAdW8uTOP24G9ABuqjcT0HDii
lT17kM6AsHbqP+kVxRfMLO6dHNIEUsEz+t2khQBPxR9w2+L6mgwVVsYy8Wg9uFSSC2JEnwB+8fBx
qi5QTIkicfTF966xHi/cYosR0yMLCbFytDEMIpP3TFS2UIgq9UE2sIlZSBPqqoPWwhA5HhEfxp9m
O9v7Z/XqK6rR2zRfBPWE9fo6DCNHblz8nSX9RLBHL+G/9e5/luY3fr8TVmLUt56tWer8w51izAjj
ib3+4et39OWuvjFzW/Pz44c4IU9UaGhZXobUozs2CYz0vZJ4H/rdw5sVEvXXCBKsF+89uIemCP69
7+0vLydZ6W20sqQJ+s9bb/BJ7lk/JcxBwsxVqdIqjTAT7WvFmyQ++Veg3eIvU83gsoVUVMww4WRk
NVh1Lm5tOUTLVPKBu1mJQLXeTUfJT2Iy0mNPDnj+Q5YtKuGitB4M3erQ6jjK2rsjzolzIl7UsZgK
Yhhm4cuCfbfZetnbPWkfJiIGpDZuCk39e5D0NJ16+QpbQDqxPPd6d2ats41PwLnaCo8M7y6nRgLu
OCaJq32Ivw2wqAFjnPHOryXsVLUtnd07E6X6s85SfOMqUGImOe+HPxhxTTX1nEXRDZztY0uNhNkx
WDQpKWp5q+06e9NYq50UoCV3bYDoAA31AA8wiUKkyOJWBMBnAPWNt8iemroQUiVeIDlU9T8pttvs
ywBdVMUS+z98Nh74QIMibqQMMdWsdi5nx80PFaPIPxkoaXPunO8HO50si74j/+gpCzEFF1nlpVYC
gutNW5H54lPN2bbcmgueAhfdLTfybgP0AKBFKqY/Rjq0WBxODd/v61OLSJkY0KYO2jXBhPIa2ubs
H2WnUbx0Eb7bgBeUJVz/RIrH1a4J9/RaGnQqFnhquo52IGKDgrDy498FY9hCHo1+si0O+Fu7XkvQ
zWPckTlyweunBHvImUJ6579xBtKkt5DoFcHsNBVQK890pJImMz2Mwk2LALB42iBvv8Xq7qHwjrvK
oDDa8O0GC/r4upl1WR7TLnYsiIWstOvhasxRdbQd4wlz5wxf0A2PtimWKHmflNPLiEydAyJ/BgCv
h5bRlCVqXHgCjy89ueWVfKJtmUbrvhma7EiEaalt6FuhhFmDYUDxmt5o2R603jyEWINBW4mKeWPM
issk4hdkTEirKdM1LytCv+RiAzCzYqj+rmm5bcXpkrLLT1lL7MQE/JusZpIx43TLzxz7gCO/RM32
aoImrLFaumBgRioml08eQUEZqiNjvOuJ6U11v9YLl3Hiut3O/EF7nrq/Sobj1BYuWohbGXk0M/Gv
V/TuJczjH8mQQIPrETweWYhxNGJ0F+EPmGWfU+R7RggJUpQBl0n0b9so3hNztnghP5F6T/90gcsB
cOY1NgnkXxT/OIjT8jiUwgLpMV6IUIh/klZhSZCTKXKvoffzOhv3h52aONhlfMafnbK44pwcHohu
wMk0SGdvYp28XKfMJb22gjrelujH4h/PYwKH0JWW0A21UNoY5XltzXw3S0WZOTNvXd8xLYsMfuPO
4u+l5IDg2FuUJoohKimHcPbuB747qbkMkR9tlVAdooGqpTOd2P4BBOIl7JXayEeXOXh+HC79XaLP
NmQddhTZgnoW35UQb+Wa4aCCzw2Z+pU7hRgDv2s8U04rEtJxGvGPBTMfXEvEGSFihjWHoNLniXEX
l9vvLHJJmnsQcuLb/YyGfO4WYuvlaT6YC/D1pEZvcpKTGgFLHUZGAHdjFm+tMAtO+UDoJRgppvSA
UhW0mOAsw97FG/5wZSbFVHb0XcN53m3xsONs13mBNzyVjcFUnRKOJvh7vQMgQAi+PzHGBa7fn+fD
pJqFSgwQdRxHGNwWfAGwF2oYfoFcFdbKZIEQoI9if3c9RwM31KClGPwHrt69Dvqh/RlGGiLagpAf
LPB3TCHBamchFddpg4HFHRUL/Nk6muAQBNY2FBmOqe4eWO2RmD716sgNPBO8tZ7cCtoKr/SQr772
OUVZeyrkP2hqZvuFOdqRK2s7KK8BvXD5eD85Rrk7K1jjobnduFqMrHyF1cytZHOl+kgKyU9yz0ox
Rhh7oycNVYYocET8E/AKCnoTgeDSepW9mjiDwiVRmN98xWBRhkW5SyrxSQCiAdrLm7GhY/MewRA0
snTVReMqWQuVxDqSCPfSHfJgGLLmvIpR0LQHKV5ay5Iz8R/8cXU2Os+0+W38qH18rjLjHEXb/9ro
zR4dn7gSo/KxGjVwUjp5Z9L/LceseRLXO3/X7v6Jbni/DUfNN4DZyGUbCpFmJnyDmKggPuXLCqWk
Ub8GWKeWCCdrLb4y6E5qyMbQ9XDmrC8XGVUt+OQNFpZlIcvDdAIs5ACUACI+FJYKy7kBlnNV8E6u
AxkCrLZ5WROWW7BIcl7nNFITGQagWGsvd+aGPwQgALsIrKVv5u6nenQUUhE1hX4igVts8qPoMCEM
bnz5ZaA4o7sBeOBNkKJ4OzB1G01PX2/7cEKnUYP10Te6lrELFhDil15Dc/R3fwMRGLmx1aD+stw6
EBtYVZbACG0Ij4CLgzPQQ2artMyhhiDnMnydY4czI/it0xKRB4z6jhzeMQxXR8TlcEqdSH6ufSg5
gZN4Ieo4B30sHctxHKCYECZ6cv1gSGARC5dAcxfzYn3bWN2maN4M9PSlQ25MJ5EqDnZkzaZOo4bQ
1BBedAFdH1toDTfNFzUll0FrkSbFdh4jOu9H1iNVMCgn1GkDQ6LwGPqFUwcM/9pzSQzeIVYZZYx8
RvsswiCKq99cyTEX+EfFC2QNc6e1WBzw+2HT9R9Zi/3risvaI2twWDeU1wi91WSozuVTI8GOMx9u
8wCUKNCjutBGSu20FDlueHmt4lKRlb7cYUCyni3FnINkkN03wvkXiD6tX8GH3eZcRuxumSXoLxuE
RoF4NkbWK4SYoEvfYM/T/SbAhee7jvOpBFJYPSSVywyxsZA/rJG0bqBNbb1JhMDXs/kECL2knS2q
lIKo98SeXg16NXoEVcpOTM8aPbwFkyl+b932PtWHuy860l5z1JzGid7kjYryCIVmStZ5S9Me/PaW
syOc/9fJPsM8oBdLK5ESOfa0L4qKz/o3xjpXLH+je07GwS90J6ESdHFmWCqVq8QP6JvnEmBAIldc
Ul5SnKu+UfUvq4mUisMacW09lTDTlRKkWWYNCxKs24A6+Oeuy2xsElHmjqTUls2JOJBE9JCkEXcx
bk3dTID/d+4Lf2RohLYO5TjQkJcFZTcob/x24G+5fub5PKl3wwx0NoxTo1b4ULgjbGElldRI3GZ1
0LzDMwh7A/kdKkcQd2ao3kri4GnzPbHvUZT81boEYtUB0gufUk3E892B0jZkpaftU30ZOgQx1LJs
/mKL0IaseoeW3GqNE9KKmwpgnTOj3L3m603wWmez3bw1rUbgctc8aOalSwNfP7qMn1d5XliMtzFb
HV29Ufyd8ZYal0mXqUOQMYJ6om1Q/pRtDXyRv+VugUT/IQSDlCWmIoRlA8BQrQfI0BecNTKhBatR
l/Frz4HVb2nahM4X8k3zoLNJgZZ+oDUVOuBg+3qoY29mTE+lpU0VHkT0pGHg3/E1pf6LVVxgwl/W
TEBCC1cEkep0sUvFfH6ukGflVrrL/2nvH9xRePvAMVyMlixhcc4t+ajk6P6TSYAoNzQAG3sGTchm
6FMM/d7786txBwwGidapboxy6NxMpblqOuG72ruAG0x/qPBMd2qAv6BpQFFnnLOgwa3d2djGXo08
RPuh6vGvQDY6LDVa4Bzj4U6PV1B4ue5F2pwSyCNodKCy6K9q4g6Rp7LGXEWESSv2KFgtgCIoGOCS
vZ8ubAlzMqIb/0F7o+TXMS2ZzUOcA/8FsDWBFPR/1WdljPlBoxUvcW8wKn7yVHdFEh0GE9hxVswk
TyhYR+VVX7r4yRK8jltZDZPMM9ZhR829CBZgBDE7/bsaO1iV2PtsUhQeO/LdkMHXa/Cx+krchTJ8
sIL/Ggf9OKQXmr9rj3IkrEX0RZ3LftyNGkf/xQnNq9GsYJHQ/hMgnTzy2SB7T+kKuEqpU+j9qwOr
10IymSwTrTweYPSo+H2o3+ON+tMq3qtvnrx0DIGrKOJO59t7uiXfYTsgm2gmkUDjk5C34DhpGhn6
nhAeyw+fBZZj0zKxTo8u7ucd0G5qTeKbirXlcdIA6rTkT+onkk7hlLnq4iu5xQ19sZpahqcdHiPw
ncP0mH8Qm0ysrF5yjEYRU9WNVIqSVu1HQ5n9NFFOh0ljWAPZ+26l6lrsflfOHC4V1oZdTRlP+cPO
c6xDsmYv4d7rqkchMIB+Ag+hM59QeW92F4qJTC9MLoiwmL8K2kBUZksHzEnN5ht3WA0AtkO4+L//
ohB8ZlNzPGuYlTxp1t4IF9WOouUnkqIFHqNem01d+r2akSgx3XQeu7d5J3XnD/JecbERXxUw/odE
cRs5vz9IDwgVnVlcHjOY3LZzZltHJMkq2ERIvoHdaodlc+LrKZ8BY8YAQdRaQYEAkyO4yc/2h/3t
uu8w2x3d5oa4kdXWUi9FNOwMTW+I8JbzFYT1l306WZh29Kar0dJDTozJoqPk6uY9FGTPAlFEhIhe
mCqmnUsfn50qtpIQ81R6q7Tgtl5yfUUKYv7w/NiQoLb7FJBGP5kn78q3G1zT84J8xkDZ+GTrorne
uXDswc4i+C0Wl9hLZRKnRYu5bbgb8Xamin2VQfUbK0WJd2DLxXdW6t59JQ9EXmZPxKKWbIZRNGBu
iv5kpNrfgpLjLTplJJ1VoGl0WIIxXm0NVkAgl1SRvzcazEgZq15LLQEY9eB36ks/sYBnwNUZXzQL
CAIwcjDNGPIS/g/bUtWbqLD6EdMovrYkSYQjko15UfmVsTn4KEbMFUa2PL61X1CadyYQb4Kiu2vg
pFb+ojBgVfLsqhuaFoJXwbTahHgkA23S5Px+asoG83wNvWkr4VWx6W6TCR54gJZqHL4C+MzyC+r0
73pU8CNPxjdLFFkKQ2f2Xoi9lzwkXal/J/wiap0N3s5YXUk1sBhO39JgKcLLqvgPPIPY08ejPesS
fubjoHkmgPRIj+Na19DtoshbYI99FeS5UAegwFfWcfL7rMc2+jo/qk1zLcsqaPmvfji92H2wDnva
k6PkDiLL2kcGTNFlO/ckks+kSvBuPQ2abxG479cJ3fivZ+whUT54j+nuxf8c0zqi6/C07EkdRZ/W
huOh8EW9w1n/7qZnhjSO8POUQFEFWzCi/oAlpc0J/vNeyGRt85miCbITxv5T2AFMrALA+hqKekIp
vmkHb1QHWf5t+4AvNQl3lib9UzWegmCkf/MFQWHOUodRcZIivb1FCEfTMI1ZXmT3M0Npvv6O5ZjC
tFd2KOQs36mJGHXDTlyiaxhx1AipwyHuqI4H9EpVqSRAOfu6nUsgwdEqGa3tlL5ks1Zs47AH/GZT
bAOGUuL7Up++oCbpSkR3E2keUWK/bKmbbH7wvimD2iU7+rzYV3ebVAcUVHhC50FAooMBXiWJBOG2
CvITnoqGWUh4FHnJUpSD9y80y7xwIwH+MR6+0rQh3TOKlTW+3zmHQjW+Sk79ESPWAV9qm/dhIOiM
pBrTpOQppvRkZ2Qajga+Cvreq1An5WYm2S66ZlOJ7u9EWFcdH8QQwI4aTiF+KpqzYK1Y1BjmSfpT
ezgT13rd81NYxm80mJxVWtYeRd4X71XRILa7MtmMBwAEmdgb3OKOMlQWTm8C4rhgs1OcqKqfOrWl
hGiEwwqdpMMMepoFJqSL9lAxGn01sMQ+mJMo1gkYZ1+VA4eI7j6gehpVT/PvkyDlZOJ4nNHInp9G
vobP6eO/0HVG94k1BkBIJmh7jnuDnJvQP46xdbx7Te6mDTkXTIm5Z+8YiaW5B8ANFeTmfaTReAwF
OxbkzgkazuOdevTuCeoEWj9A0cXdiibgRGw0NgHYUPC9wK1sX3kzCo8GVAnGytF8lx1JhOaCGg1K
it1vYZMUAI5lzlfGyF6QsTjZI7jrNY6/rMPnkCaC1Nuj6+r0xvEuWrFGUPGFFpW3ogHRsekAepiB
qOvrxoRuBh/4JVhbGlqs94Sz//RXiZSO3rzJttDpMbnPwVSsLa/MgpsnK09Uz5Y8vqHjzCymcV/H
yhIDs6qOSPwRDAyGjKoYQCPNEYvZtHfFNb5V69eItZxTO0fz5IlRdMN90OuonFe8F844b7PcZ+F/
zMt+FZWSQ1cjGkZxpXEA0FER0Aqr3196cn7K8SDXCptxrM/6wIWYjlKf6ww6Yq2BjDlClsnvH3kp
qAOBiqZe3OOwfJnOVTrBYTaUUi7oNSrAmvsIM88WDB0lLKamj0aAod1I6h+mllXOl7JPi48fmZlE
PVkm/PlN1uuk9A7kn5HwQAzYkEIPl4UZBriLVlT3ZCHx4zZSINAwSgcKy2/VdRnVr+sEafOC/GGg
rrkDs2wXQlCO1Nmi6Y+HNaFV4vUqv8OWGtJpqvcLi1oNE+GruyKzn9QWgx1YSItLa2xyDHFGGOrg
zAVIk2lZhzRcVfMMuw/3H2KqGr1IlAisM36Mdww91gI3u3PSrAUmHPci8zZco/6ewTTL9SIfC/yW
EmcKPLi/PqIwX1h+88qh0h78e23l6EgaZB43d6wHZ/2EMC0dZsgJAh0/+8fEfOrrZfLb/tj0nBN4
LEHsXpO1lG9G2SfplruGApQo4jCGJpuspXXn12r7E41xQBqAOHunJLcSeBJ5fr4nWoOXPFJsS2De
n4PPXYWDMXx7M/oE1RwtWZ2MxT2AFxI7yw6W8lhbChQnJATRLCBRw2VdJ24kzFLFFi9y2jl401PE
aCVtqxZwxzd154n/+eO/t1VzWQpE4KzDjZqEj8HtvNdn9cnKp8HqLDfb6b22as5r1CZtOe8qE0bC
e16525ImwMMALhqmoTPAqWGiSDztj9ZKgVaXzLY8szoXl7yhPrUif2yHhv5mEkBF/Y3Mt2xfGKbd
grmUIabjym+8Whz/1GJOb1XCSIG/Tdr8jNAl6sIe2Y/Kq4dhLE/vm/Uxe+tJwTyDSbWf30mR8G3v
E3jPpsicEW749oD/CWYlgJj8tT/WE9w+xYfHZkcbxrWNWIXpkiUfsru76Kj0NPZQbULPH6XYowGz
TPZw5/cYUTGVWlAqZGyD1WhfNSkkmrdLTvCmkZTNASfmiI2Nop3W2Ge+Y9EcFKREjwCNYpWKBaa2
bZ6aQVUehjeshD8XhGO0HERSc+CXWH3Cez+6M2S+2FhjrIA4NIQTT54MMmUUQ0VKXzdiBn1HZYFF
0NYAfCOdFFPpeVyn5CZF1nBmLzqIjezVliVf776zcHbghYZMchwhvx8finSImqXSA7xX/vdrirnu
qD5oOfzjiptTsz3DZWcsiFqkurq4gtUCCOWEYl1n8RNxv2sW+asKyilhqB6nPezJlxYNDoHn8BCC
l0FCTpsWVZ8j/2quS0uRRFn0fX6yxcv/BFhWWmbYpLGTgVkO0sBDZh3nSQxBTFZeYzstJkxmcMm7
u++FkUZ46QifuNIEKxLkM0oOgGpQFctqoV/+1x8aIFiAmfJaRTJetlKC+tBEYJ782NqT0G1qlSe0
jVHFXvgubhs98n/abTFanaoZpDDLBilwRAeiMosfjQhonxn03yn//1eWr9THS78oFdPRw0bpw5wu
DjrxGHG/rGB2eHxhvuziSktElJ2cdTU4Pf74Lg+N9jn3PYwxelAzzj8uUhiK+gF2j33LMvTF9W0Z
oujD8oJL/OBAeN1FeGdMuVjkGpAcISD4OQRVX/3ic9RNFVQwIqp3v57qDjdvplIdMucSNq/4/qtw
svqX5IbfGcl+dFER4lA7nOJPVlmz4KRxLRMpm6ZOFM4h1MFtX4REwaZu2OQ+Wn8TqPoj9bIHsYns
h+PwYEC+IjeuUjqf/FSqpouLoNNy+Z9kXgYawHF9g5r9f1v+dD+1rkDM6DykSLUWTPB+g/dk71gX
tb36H9ZUjM2TYG7kT4xJrrdbTc0jVQkmxhHlN/Jfk5cty+GI+/ElNkD3SMoPlxf1EyQoH4+OO/K+
Is75tm5gM4TMWOnIOLI3J2O3DbDMcCpTJPfLRxBl1o+z9MK8nIn/Vrzw2ubIEOlMBLyFzpAw4hqu
cPY4wgjgTfcYKOgGdmDiqOW3Y8yv6gELZHhdeS6MyCO/uy3mmEm+ypLaBi5ZOQI0uZerwAug0geI
46evpB/zUaMcvj1aEe7wLOYhRQQFIcbrcAepTbo2Odajq3sf8cOQiwJuYfnOvupqsCn5WT5fKNv7
8+/5zihfO9ZuAC+FBbcCJOHmT8rPjU1ZYFxTq7C1W6PesiodxsXo6tt5VsOYeMs7xtgRNmXEe3hJ
gNWGurrSY+uoqmJhWnenobjbciysBlA4q3kvhuzpBdFq6DDTsczwZwOCDBrMFf7fgpxD9TIC4UeH
+HG0YIydE/mXrOj7FZ2XGIbbmO2eC1k53EShlKc8tkWgC9HsIYm7P/vzF4wGyF02SMNNZjksy3Ji
k8ABicKPg3z0pSpMwo/piKcyMyn38O1aLzNB+9VY2G0JKqBLuu+/GetdHx/QZustiA3Gz5R15/z6
JSbfO73Lyb2DRRqZuhqNAeN5CYysdWSWE1nFipHbd2W7OzPSpU3xmbV/P/HNMjppwk0XHb4Xc6Fr
8RiOFeItdq22yjOLIVTT+AHPbZRc3UfraIUNFsEie+FgOt76ceOJUU68X0Y1tNUC/t1ilEZm+mWJ
DOuFWYPF5B9EwHJWatPL+S1PbPsbsMT6hBsnDPJMEI0Wbt9hUVkNu3pE6HM7MeJ4ALEdbpfFejCC
4aXRNa1mF2kzE8o9Y/2Kudq1SpvL3ElX6HeHPKsDv+ccS/eet3ZVME6Fz3Vm/1Eh9qD1ZNr8IwwU
1VVHNoXhUqVMsaAr/LMrSsueaG3uYHMYeZj1BeOSK5anf8VxSpI07qozHXg6IUqFWqIyV6f+dZYq
x08j8A2rFk8nyo2/vEDzPry9A+eBsYxT1HjV6kTmHJlJAbsEr4Nw74nYNUr7j1hWtukouYelbvfq
ZxKPc7UB3PoeJM5w73ndVss0wlNTay9N9DzHAWIe7Z5R3lp29qb6Keb6UOZiWXrtN0vK0ZQginIt
IIHWtR6SJ61irIdDbfz3nay16F5Es21rTjZF5BtI6PtvcYhRMNgUQdgIGUbdGRC+O0cwpiFeTBJK
yqgdZnOVn91tEFrgF98xyn5M7r/XaZ7LSfhxh1MJMAdPAy99laxMEOrAdfskHMxOcyusIeuXWEXQ
DKW6/pCpxy4pryAJOkrXsVMsR0i8NF0QFRq1KUXtwpLQiX9pgifGvinH86OPbTZLJ2wIA8DKkZ8B
hpZyAFeZbmjIAlRb+AgHevETOSf0naQPlIsPFAi5zsSP/nq+a9cYdvFLxSR0zYigV6X8EMk4O0hJ
Q3kYu0oyVLgQ9JC/mm529OoFpyrtpOyM0mFSbO7CSduU7eQpUQZMiT5QVjVTs7CkdSxyI5/QlrCj
Xt806IeARYYEXA4W2HEi+B5HUr+LeeDLgWa4Bpozf6uht6Z64/FUSds9EgZRV0bpliRMLlcOzueC
i5IZdnxKe3c4WxrFQiFCOXiq/yCCsiasAwqTbL5Y+hJNyIIQHgNImEpPRIaYQE99KyGxFymCHcFr
xOqs0snrrf0iJYO5FZ1glttwy9Y2yN+I8iy34hFKdiXCZnISudeE+fWxV4TPJeCO+/p8hO+aOEPD
AqFCfa10Z8T/0QIos9giEQfBun0IfuzzSZ+JEBsdu1NU/XsIFK/NK8jbZE9ouzQJSc2mBwUWiCU8
HSDo27ROw/02hIyLy+jg1Uefribkd71pwUtlgXrdC7p+02xa0GgixSlDh3ZYtsnhsjbkurpVs4M+
ikX7YRSFevy5kx/+D8OPVpq89Ej+Y1z9VWDIbq2zexf+wVC9MCjGUdI3SNFxYQmcylLjJe/Fzw1m
gZDkROEmWQ/X/B+N5Ha7NdcuCTPFJjZJsJMFqQ3+Ib+mY501yf/scdyzmmMhk6f1TNoHG8jtJQ0j
KPCz2YEO5gG2ybYHrFOaEhHKShoj2W2J6+MTeWu+UVxl0y+wLBeMA4LwgN3bN9WNet5j2awrHbQv
T8WxD4SdIFMJMK9ixc+xZP46imAQYUTz8zyptZoYOZdKmr9iluIgk8nYUWfP0yvYxiWKsb5egGnQ
FSYaUq8pWS/Ql4m4wRj+S6tJooxhyS4TmbH/YYKSx3AZx8NktYnYj3+DjUgC2A5TGQToQaPvKrWU
UmhBOABAGTagNi2Ih/prbePNNTv5HewAgDdke6MkkOatsk4PRLxs8iDo57YOXiYKiTQ5g3bwuryY
5RV/zpd0QciRH/rlINY5aXoFPMNlrsz3NEWRPRs0bEs0D8wDQeotUAcW17wvtVGepkgKro1MNBBa
T1fnuL5j14WUinMi05GxMnbITI0x3zbVagqhTRkEtWfVvzhkA++8hLiAi2a+YatRRRQuz2Ojt/6L
7EHy71HE+J8a4onZ3HNj3clNs0s053hM/FsSipHVISMxGv7F5XYl38ZJiVkrAdbamCVd0CtnrRWI
XH+uQGi339x9Y00B5v+eiJ3k3gb/RAXHtQYce2/Bk3rlM6NIl4uhfUSAGiv9+XIYOYouBA6sB5Sb
GFq+zMeA1qyeTusEunJydNAHfThMUuvm317JLwQpL8ijs6GZ8TEya9aPBzJe2t01tERA7lJmtg8c
5zEpxQ/7SXGW5FHzDQOuUaNQReqDf0D+nGR0/1147CcmlVrp6O/Vl2iO4Ro17ByYLvQGOK7+OFLf
QZNLxZqWBTo3GbdzHEawcspfJM2wtTfdX6ofcvH0Nk9m31iY1+ET2ACUVhLwF5xTpOHcdWs0CNgn
hfZx/ZchwUuujxias1jfYpS8pjQBHcnDyvUKeK3hJ/2goPRhBiCSqoTJoSjXXUhS1CR60wwsidcs
L2WhtYxW34PtV4MJsU/ZHBtq4C7/SuvmGi8ud+xxo3eGpHq32Q45mXRamxwG30r6OsL4fvKHXm6E
304aCUaz2hM0+ONwFheq6pnCuop6eb8IuveSkcdhGqUFHt7gq7yzcPVkRtLn01MYrRttTDNwoZ7N
V36eotWzr4t8TB3Y7KcRJ93+CPJu7C7lpt79QeLYiCWuPmxQHtu1xXYQZ76A567mFtRp+VGzgETi
G4XFsq9FaSdgm5L5sUhFj5dwo2y7trNfnjzZfH2ojTRYkUai6FL3SqcaWiNhzIj0Fgyiq1EVoiPz
waTsyWb8/wWMJK1//2Ro7csjcH0fonV4gtR6VaRXgXRzlL92G7DV1jKmUbVT4VHoeTJKXrp3/9KT
4PFdQyCT+jh5dsWxMJZkmyvlgCgT+kVfrlC3QnxM4NM+3KkqpXvFHlhgsrMgblojAIgXBdr/1+vk
FoehTb3G/nlYn2fz/TIS+CyUZCjAtzWQk2orxlwvj6I7xLrYM3RSNGxvEPQgWkDucmFqANN3ovbJ
wXnLHlDWYL+cWAr6ugU6ix6cYLiWldde/DRAbfFXV5dgR4oXg+Nkac0ET3rb9udg2hOAaUss+q7G
ExzvBenA38L4wkeksBmheq2nvLn9fqmdpKv2y6JDdmKTFdqEbcwg4xQXFoChyODxj0xIMfgUluv0
1H8b9y9cL6otR5MMGh0XfkXujt8Rri9p91I7miTw1o69lOkx6VpjURWATMi7cs3B5B7zGbdVVg6K
9YqOdz6zAU4euErVHclJnZ201t4y45sChLFxFiewFI4bBiFzx8BhrcLrgO3vrC8O0kdLxItEJMEM
sKSyp0hqA9oXwGPu801S0HIHYFepQcv6Zpnp8w62eE7vAp6UQ208Lg3xm3irRdfTsrB3K+DcX/Vt
fKCMAW1mQvcCfZ9vdN7AYtzIuDcY8cOQk2Sr3btZs8WNZw66rsrtfoSRBMx+3M3gPIVgdjkE1U1z
S24NJPIStCQyAhqlj6UMGr8DyYMQj5ON/uS5e9HnRAaQ//x4/VE2IN3CuriMazji9rO8L3n8Zk8q
cVx/Xrahug+MSQ0++zNb6DGV1lkOb0xaLctGbD486xeH7dyjpENYUYZFD6ldNwTmMON5R1PZ+TXn
MO6dJLvwmAmCzW/a5UbNcm9tpuNPZDXO+/UV7vCWMiIiGORHbK9z19pUX2fHPfObfgweORAir1NJ
0KZpUzWgHJRwOJNF1bfkZIFyMP/3KNRk0wjqmxsSWX16D5mj7exqHlr4Baa//ZBfNnJ2MKHmNUty
cCFb5VvvXldMKj2GIrnkFX9qNIdtTIZVptwyUF5KGbeblGkuIEhWZsWR6uTLrIavFRJVcPPa+rqG
kugi/IyVkmnoLxjx6hMr5WD0Hp+wDzYn13moyc5SyN+vFw+cv4i83iGGdwtnyRsS/6fuuiqpZ9wA
BzZNLr6/WDCzL8zangrtwtHFqAyqLn4dWaTuJ8ZLSiAnFN/onzab9lY7XHZKaABLpa5uHh1d4dkv
INK3tX7En7pwDrFpww4o342Mn6Yg/r7XXb0Us98WrFisULpVhO3aEcTH/bPfg+8WfsA+QHHzD0bH
NxH5TQrpphafOGUHPOQIRIlV3sksxAAzqFrShElmBb60R5H4TKYxMeKuAE2CgHx58DIjwjqJCrUZ
5hJs/+rZ5vQ4pogABBP6cQ92AfQANy+2PgJB6aWYzQCtPpLOYnyELKaNLY+5Ye7HAYHNd6hzg5H8
mqrB/GhzKMWPD0LOnZY83jYmN+xz3Lwq/Tc8GN3xqGl+IflQ6sPLKbfFbSpSXm64+5WFauSPA9vF
1VV6ELmgKaoULdTZ/x9+Inej8SovA24qin9UodSBThKvMuEiWNngb/GbBt6WTvp3x/vzlCDSbd7f
mTGSrcZAoreYSrKGBIw4s9+xmap4PsP2z6vjlLPn/oK80nz+WEdb6oTbTiOGcEJ+fdVfQmxTVcl1
ZN1rpJ1P2iUJnVLMLTXGsF0qHlB0AgGczjf0MaZ5Cafi/6o7ecfyqIFVAWt6b98r89gYM0oto5F1
h2SFo6HSf5FUUm8XXz+OUXLuqN/XfkzHNDZEqSO+x6Hgj2v08Yl26aTGxZyloremWhS8VDnOiJI3
5NcVdKRtFjeDmwB9/veLJorEfuUejy88ShptSpiSjuIJt8mwEeODqZBZz4bk9gdjyvyNYAuhjuDG
fri/UbBb4ht+pVZKudDA6NMpPKoJrm0CJjCylWfzHBtmV1yIUx9ChffK6tn6CFZN5KOPPCe6kiK8
vNanTBcJJlH822hsDeDUI3DyTinS1yfjxU9N41LFyQUZ+fQXiDv0A4K/sFEZ/caej37BeBhrg9Zm
ofxws/H08xKdwnDaioKjS2c/Wiof5ldQ8OW+lbXNJszY8VFyb22sTvba70PFlRbGivwKFo7OhIl6
klaqJWRF+yOWCUQ28lBmi2beL5KeIOkpulXpu+LUFfA+gOPR/TuwrvqTq5wakw2s73g75ARDAB2Z
yfUka4GAPla1amiwPcIhY9A+Fmy0Vn80fNOOLsivaXSeICfYE7lDQ3yX+YqaHvADuRhYOrVd6EsT
+LabKSUpKjN54ZEMOa/+oTNG3aBHxGNZwCSuCfe52j+0x+NrY+d8k/R9/4mxDgGgxaBfzEW65A7o
bX6XGCi43j8SAKcBktSw0phhQNBlzgTjE9cXbb4+XARQQ4mePtsSVbAajY1LiejnBIYDIvH5l2/v
9EPD2nU0N2MlQRrQ7jTkb/DCjwvg+ofWpzbSGUc5S4e+TJ8EY9hK6IMrAbDPIr+E1lOZMQMZ0/Vv
r9e97YFlqRvpOICx3jhQ45fOpqMmO4H3m355jYecrjwiGex0+qKPQmq/FRRd7jI2Qv7y98fe+8u+
LSGZlh/dLvhPuHGD1sZ38QbVLbirm1hTX1PL3gQ265yrUGI2FNf35IJnEoF6aXDR97Bao4En479Q
WcX6fU13PASnjFbyzCz47XqOFO49N3CvBJt13Mur3+keeszwl8Iq6uiH0XyZO/fFt81ua2L1Qr4P
1f7rh5VrAl+w2hbDDVBEgorgpEzGkow2jt8UrtP/gtdoMq9avuVWapCfBAqj9LsCOUYQnsj/55Ck
EY2m/Iw22KiHtNJWmXm5T7EGl58CPHb1I+dpKiiGvE8ecb1TxX9Q4Ji7JTw0OKsTy1LY54O+3xXd
CcCY4so+ShZEqt2l28BBWyoesLIj3XeNMwbCHgLNwVhXy7QmEGG8FfRyQjglsD44YpGTTKFJ9vAE
QoNZJSAZjGT1RR5PehEtuisZAMOm3oj8LFHhk+zfegpctIfy3Qbswei6uwbNlk418hBlCBDs4Qo2
SodXx7omWGtk/OQTs8OnSMI7s08qJipN2nR5nzyYcw7mSUc8Fh0iuSq8WhR6P16KEl164GFg7ZgQ
3vzcr/sGYI5T4DbWWyqetoR5uyntUfcG1VnW8gr1veN+b/onGfMMQs6h8YNlvXLix0hLrmTPyyrl
gLf+qSMPn6YbndSZERLGzVugPM5TpDn+UIS7MEIy0nuObTE9lBzLaOuaM/JT3tBHmgglp8f0b2Rz
P5W5JF9rz/i40HP81h1d8gjVxbRDbkym3cHzgZOvJ3f5nTmg4o1o5E8jyl53iL3g6ebyFUhfoCu8
MIkNfAQl5WrqSQzOypzaKxtWaFsCrzHDt0lELRjnFWlMvgOdZfE25cjsekE3tzHoLCk1vj8KJEKF
8pFJBSFTMnCX64kVZllK4OeD8qA0sMIVvslAdHHWHvoUuS1yvPnC2w+J6IoaL+Cc3msoCDjoYoZC
4kbMebzjVPQ2YJ0W8OwZlmh92IuWxav4guOKHX1xNA8ciOZpyGE/Z0A/83GVUoGIeyBrEaZbgLBF
+52sBpcyzb883GosfJ/jP5b08qV3bav+ILZBAIlPr5hRdjUBKJLgDgv6D90NhMNxsIwwJ+vw4ppT
e3bg4pwt4KZqPjGKPfzl7Hd0JskleJ9fyp0Rp/N2qBkKrQz0vTl4Mf38tVVt5IX4NJuKVUeTwRyk
09Ce+DFGUd+FHPwOm9gyFDBm4RIloAgf0rQR9NE0taKAS2suE+mZDJjCy1P9NyVeAXAIOTuhriVL
0zHVWsBkCuy/1ZfH37Wc7b1eiKfgLtGdvc2FmRnsv9Tz6g+pJA23Rrua4lnPevFUaY3SMuAfvA3S
mvTC9z1rdY3nxuEvQpA7PCxlB2CuZenh3LNzowOBsLUk/xj6kHtb9poXWrNkuP/j90TNNl7lg7lj
hNuuu3fw54tRB4ch28C42uV0qj0psosO7dAROTbeMsubmkiMRiTJtYUFYRdlDOjOOcuFiOqjwkB2
mgxiMOBlkLt3eGDIyD/iZRcZyZIf2VCG8eLNzMWaZJ1S5CUg50AB77Op4eJNqrIS5SF3XqoWcqiM
2qWJKdk/jrYb6MpNXrpwV8LYAzW/sL18Z6zL/Oa63P2p6hJlYjZD+ttEhPB9fkia6JKhVPZ5jQYd
rsAQFqGiklUDQaRD+zXnh02Ow8DO3uV2Xu5qbJJ9KYblMs5eE+PSVFEa4SWJBKjffmg8Ypd1DLc5
h0ubB4DGJsgGPFBpGGytFnjHsFNzd6dj00zpGGnTPRXwFCpdswLtyAo17J80IDSdoQRSQ/F+wfXK
5+69drJ8Spvj99U2eY9pg6hfZGTc46qbt5hPLZkcJ22ffaBdqZgBidQMWlkpVHSH0UCohJZ4fTNV
qe2+xysynijEv7vO03GplJhPq2MryhzSRqTkHYn78fo5PUhsK027nYReQsvg0HSqaBpswEAFDuHx
H6RVDCvIez5nlnkL256OTAsvhJ45Kx1T7rJO/GQGSxmU9xMcl17wfAJyFookR0Db8LuuOR9oFv2B
Bky9hsjVREr0Klpoi/FBxxdIV75iaJ0AY6x9hNX4VmitJ3TrvTLnQDzwqXhaiZdqbzn/ak7qZe8A
YdymAF/iCLeIm7Pz+AKxpCTJ07idp6pDqPG5r8gaYmVoLHEaHCj1epZ8/aBlqvIH+5S2IR2cob1T
i6ZeiiKqJhQoH7qoNlfU15fOPtf1jsLYSsr9AIppQDBfcv2bqEGrdZlgYcC1qA+lBe46C0Mrlw89
cpu/Ndzvj8DYoXQvxLtnRUw1/hElSHY60QpD8dTclJdWSFbAHAgIc+AkftVmi01MFT5J4tOk6BSt
COdwTyCkDYv8U7zvEBtX5wFthfclkQJf+PTlUfXkr2JGQd1f5KsFwzfoVoLlTVXI2ocVnCqxk9PU
JK0LrcB4u0D0DnQg9dT2QTk7GpDDetdwOMvVTmd7CYvBGNw9zgkwlCMaQeWWzHxUlYn0oX7gV66y
yF+CauEik1KcblRX8amserARCos62BZRyzYFLFSxCD9Ox2PbauOL4M2nhyK4DIZiTZ8vpLlUleCN
7UyrbnTRUYVR1TAkR/OJvOXcA+yGbeXPTOJKetw3A39o+pUvyS6/Cor1Y09koPT0sLdVMV0WvL1B
6BiYmynwNZrEU90zXGhsJ00uigSV1OIATku5/3sE1UkeCnZvzr+gB0KTFbev0Prgb6J6RZ96+/bP
PMruQ1QNZk+7QCGbwvBvfdjt+mRjGS6YrzcWTx9Je40Sf6Q86CSLR+ABJ/v9PAobzOeFZE1lodFU
PwsyC6ytAu1UEzvvW1N+ooFWtHTIVnOU6gPiD1oaybEI54fqJUSWFc28qP1CJ/1YyFloqxGlwCsQ
c7gGF0WtCgvEnALFfWXAmfuo3XX3ZNmjYFPIwg0D1UuMc1XNJnnBArlSva9mRpLJ7FjaI7R0D+Zm
bPbKiLXeX7eZKM+aE+sMEzGelDzDFL0BbBOJRwANbA8VGXTO3U3/oBTsfbViEJMw3FJNMdADNEoc
yw0ziiLZr2OSqWraE1Km57NQw52u+ObBn/Ikae11dJfsvacjO0IyoSYSBqrMbg5U1qRMAkE3uoFc
RcgsLfqJUmHi+eUUlxBQmDIRi4HPg3SUfg+qxX5p2VZrH8sIdR9lgH9iuLM5NgktqmhNE7/ga2O7
XPj+qmGId5GU3hJ+LwB+tA2CIkp1FI4++16Weuedsvf/Z6lmjizECGGrB8R9fDeKsuDrnAbS/X1Q
fDFtI+OhEEzYVnxEGTNgUTwK0Z/d2xKc9UBtpNVS23ZxqTHE1m7WKZMASSaXKHrNfsTAIuxSEW9i
hMhml8SGHN9dSN6x5EQRWvPzc96EMKJBYa4cyCMXKUogb9oa4ikXR+e+9W0F7gVcLiWbLJ9foCdB
Jm6PYWNgdxzOXO7kARDOpUEN8765LjQ7VqNl8CXSjRNkPxw+110Q4V5ersb0DZczFzB+dhx4qZoU
zDaN/xBp+EWTYqDErqYW2N/InS/BnCdtJa1SmRP45KAhZnZVScY+7zrFGIBBFA1zqi6OoGXAuSpc
d3Xmo1fsa3/rBaCU63Q5reFK5qhcsbIKO8cIGx+Jee/jfF4U/YPiMWNEznBl5rJqRv3NiGN0F2sG
h8fVSUQQCoPU5l+xVHX5pwnexSFuivDYQ/Xsn90VqRrSixLiA7AZ1lB/5lLclcmuMXqX5GVjhTDK
s/Gej4iQ35afYxDkjY5vgG9324XoGMzJsQ4FIVnC+OEsOak24e78Az2aVGpuMtENom3eimBhRJVV
okiL2bRJ70Qi0GeSquzaBVLclR29C/fd+9QtTDY/wOXd318qgY363HOQA6oWm01xgSnYFzMinRiw
VLpsTrdnGl1KNnUnmMWmex0VILb7s4Tuqv8NUk6Gr13NzvrjwhhIQIuueyi1VsOso6BNHjN6jNm0
oUZ3/KjCz6CgyOoOmwBx1z4VpMTu6tsEM40JuTNl3LC6Xk9NO7qVYXQnv743wSmt/LIGcYijTXPr
HhzfXUt/fsOnyc335IOmqvoYqD67cemWPjpwKOksU5z6GGmSIuGOHv3ZY3yR1S0gzLk4X4hzMEKV
EZCFIfCvly3GY0FQnOa4E6XXp0/PSOd6AEYWro1wa7AGUvCvLI5h2o+fWMBUdzZoBfe2W7bcHdf4
a2UP3sA0AL+SVmmWXtCGEf6kW1yAHTG7OR+86Cjd7UHVnq+Xwqei3vVTsRnY0agnHyATz8pvJ829
G9BnowvFwrKFejgG/QPwR3kONi2GLP5LmLa0jeSO3liqrJersIzHiRzaJCfm3dRhtWWo5Z46fJ3W
4+KOa48jJjFc2tW8DNHTeB1B2hE6l1dF9l3UCw3o1kUPKI/IoepXf7jseAgN1OZ9jlXwNiVYnEwZ
xVGBlMyDJ/PJI820jNBqrvsp5XhQUzjNj38VArB7Zo/P9duz8yVAdcbP4D9YGPuc1kiiV/4bG9rR
FDmPjT7Vkvf0ujZo03wuGJYnNWB6O/hjBvAPlVg+VjO16UoO3bkCZHimyMUxHrb3kuy6l2Zj2vPm
MhSzyUx59GqnZnHwtosBi8FxiWn7phXdSDah5SQtNK9+MTtG7ffLMOrMbMyBmyY8Wplw6u0kKSLX
8Ss11Eeo0KgVs8/03JOyx/nXqny2JHR8w/sP+ZMR22LFzbCE+OOgvxl4yquOvKqa4vu/vqK7csTN
b+dL+20eJtPZYgaF0Z5pAgTJMu7c6X1l1ihD0ks7MiQlJ6DOIJE5oRSEKmizAFPPGQtdSEsj7tYm
oYw6KQRhC0O7lbhyzQNBRDmIUoIavcSKePR4DfXEfOqv+/3CT+2Qo1paAXR7+3/u10QES0cNYXTR
PfQZaT/EOm0Ad9sbscFgIUZZIA/j+mH7nkzIBxxpovaYJx2eYkezQKDNgCVW6/3RXhP6ioBquhD+
jLT83LO0mkFhzsXWaQw3a5kscGe5IvgC/Q/egkZhlKLF6q3xAoA8ToLbwfLug4n0bENBKLj1BBNf
9iC2T/NpnJNSvZsaF0PuVojPc9e7xina1RSu1w1OK/FrTQbzAV93Zpib+zTWrHFHWonQqZlAqQM/
0bp9EnmTfkQiYpOeNlt30JEixSRYXK1s9IofVDSF9ogjeIJQMaPWs1xHwkwaZLhlpq0naipHM8mv
zIJrKrzhbL3NTkH3bTet7b4Ld/SK3X4H29Goj+G8v5QzW5RltgOc5/S4H9XQyOuArWATIKki0ksG
yMHelW6DbyYer1zxB0UAk0uIweG147SGR1M28gqWtXwGbP/qWdDt5UhUJ7JF4S4Af47w0ozrRhJ6
L12Xna71h9MSUzQCdMlOWEJ9bXley2EeYuOgZpKr5vdEqo45pnaCc2qpwKStbyxArQdDpoRJVdeo
E1Nn7vxHOMQPBbwxh8eViiazlYxhMTLAp4gQtY5Bjx+qKoLEj8UMycrQStJsFN36BPXzKZPW1WGI
Xs96GrpTdbHcdps78KkeiBnjvdtBXr96QbwRfwciU+7yq9SX+QY4k1cRHZNUTcFLtnNvsKRjhS0k
QCzeDFrDRsJB/7rYJqRJLynD7Xn/J70Od5ZuoekgXrWZk7Yi/4hXgWU3hvfBbUiChuzBFCsfbBhj
5PzWCdCMVV81UEAakit5RBwOJYnVX2Y+STV2gT2jt4nWulMRyb072PsSjTauCtKN32HjO95ZsuA8
nohQir3HnFWdJ28oxGcDhHPmpBjlKm+d6We8H1arVkDJLwfrDdFBRG43N3Ew6Icwlbq5msdELX5L
xLtU4WelBXjAxD8cx4yGbXJunfnPTqZlcl/XDi3YRabny+sIal1y1n55/hHiU5n+mxTr5GJxI8wK
qM1XZ5jZy+M+kNz2TKJnOnhoXeJOLGyV1SQXYUnYKxIC/kOUp6U993jXllCaPoPilo3THOtWdiKf
VLNmqKKaAl9+Ke6Zy6bCTTbws/OdgiYR2kvB9gViQT5feyiR0pl1glImp1rgYYuf9bj80ANg2UoX
vT8dMdNpD1uyXXWeSIQh/ojFFFXtccuhwRVGjsMvfb8GneRo07Sv7xEMM+vtWFW9rp8PkxIwIMOh
6h4D+a6BnibDOgRIfp6aoXtUz2TVQkn5lBOUDUpx76ScFgKkTQe6L4ilWLh26Jm4AmLx6MOEXfE5
uc39SFBEk42QT0hNLdBsgjR6NEsp3k7mXZRiZQLIUGtIhRNchpqAQijw8e9R6H857jPSVbJ+Dw/H
+S6vWevXt9cwFyXzTVL6r6wngB5DOnA961qECoGCn8DG1ZS0EfcCCh+LQ+4hyT8sG7I8tJz8Ayb6
IvNkIOCh2d5avcpJ3XHdPAuYd5DwqvbpPQWI1vus7PJ15Yn2U+EECPl+N0ZhKSF7vKVvgYYdhPt/
WI2xBIR59mrUG7pCWGlOwczxtSlGV7tgW7uKGhRyz9dDT5BGQJ4NiQYvuZuUH0lGaCuM2fOm4MvH
uRHSsl4AkLoyWGarFiDDlbTxYE5gi1GO5byNHAN3T8XFBBjRJARuLC73dn0dFSv2MUs3BKOTbV4/
Kn01DTbdj1rWPZi7bKqLYK5ghijO+krirEarIFJddY8h6UeuZMI/2IhKCKXv8Jfwy12tJgADxK3q
FviJpKsf93f0otSExIgwgmCFuE4p4xbbtMj/feChWmTMkYcrGXQlu2mzGnF7U1OyP3v+uUncRrNo
Or/T1CIfnoX9mWbY49o41i5s0fEIutcsGC9bhmRqsTIgl8MklCGB3USJOBtmzopI5JFvvoJ14U7p
AqxakkYZ12uTXwBQkNHdX+s629uTdQp5q+AnC3Gbnyyr8MeuZam+LTTT9Bf7yorWxYXiSRp66XjN
D5i69Qd13hieNeO8jTOXSyG/zQmGPi9bitH2kG945NrDVbmfXjMiKh8Gn9wHdRe2PLbu0gxpotUV
mq+BBmvkcKL9Zt6fQKmmVCN60yrPM2Tv4o/TaM+AD4DFiKfavD6gtFM0e3etHXlzEHpSv78JCTU3
45dWrHhXZeAFbEOi/5qenEBsidj7UVWGlxm8vtyu7AQbvUNyF2f0WnfiCmIZa3dTSZtJGMBABn6+
Rpv9i9k8RyYC16MlcWtgmsPrgrkQbPSfRrlanVmHFYJGlaVStK7cXJzANj29WNx+FzCpA1lWeUQj
bNjjku/DEqSQ6VPSQmp/L7KKvabZJQBp/DN/U+PWtdKu67wOP4Zm4RufqR3oGF3ZmhDbhX0Ocnrt
rRfiTkjwDz/JsBd0OG1EFGZbn7Bpv54ZkfkvR0mbjGGPLzMWBsPheUDO7nblZP2xCSgqoTx4ieLn
mJHedS2yfcJvD8nVzVM1y4ctdnl9HtO7ZOFeginfIPjIgbG4AbDfwbe0fhVuqp4God61g21sbIin
xFm+sKCrpwkVmPaKx0mW2J2euz21bY94I30pq6Up+t5WIXy65dxylsOx6qu+fF9bP43py8MAxANh
AeJAGBEt8rnwVynCB+WAzq+JlRUI6j56ARhWYwpLcFl6gH8QF+XU9QAi/5WvNqPg66wb2vL1arK5
VR37Pe/WuuZd5i2hdyiIk4TZ+P1oL4PrfL8FtftzZ2xWNvwJ4CYHBJl+F0Nk6oxj0s0HsoS5F+no
jCdv98/X5BnvRJNdNUnHt2ZRXe4pWxgep4ly9yx/KWjfFAUArWHMVOLOQXjM7ULPVizP5BxwemZ8
97Li3KNWuFtsShKuKbLpKDw2BRT+rXoguLIwRsQlPg4HXwYCR6gVif7gtWTPUWN2FgZ5TOz2HWjO
Ilt5mx8JnfCZpZBOAuL6+RQBf97xzmGwa/kOt5JBhV2limF1wqpfMsSw4VzvnysNGictksxWf+Mb
PC5lHcT5z36DpKH9ogYSV9R75uUHR9e+PBbjCopCwBNgvQkPQ4Ru4ttNpIU9LYBuuVBtPzIfsaOZ
xWv50L6bYsphSLjwW4WqCIQZXzlGsHBzQ7U7drpASOlhEy/WVbLgQCpsWvMiaHYuQ+38Yhdos78B
rhs6+/Qu9/pvbPUu7rQepI+CNj/csuwQm7O25oFistp3z26VePpZlzqDKlkpMpi60LuJ3ePjFpZC
0zEyjPYs+lR4wLGNfvdjfaaDpHecDsSv7rJKjoSnNFFZ4EPU79Qpx+VpIwxqRcSCVnZMQUog888m
vV98PpkwkJh/36jXbh4PT/Bd7/Q7RmgFCmmQ3CzIIukjwUi0I8+VKWOjcgEhWpXKW9EPtC1wdEvd
HtOin+0VCDooxJOv6V/F/aQTK4f7wL1KP2pIkx9KQsIndL6wB0o2iRPW7/IwGDZ+YPYqWNkK8Pi1
Dnn/mbNcVhEp8pUVS4B5+Gh2+aUyDgEBxe3ZV25q5ldTKovBpKqUI0DfeBVJOLguaekN+GGi9tSM
lJ8jCqJO8nco2DafPoXol7A/82VbkD15EGLPdsxDnf75Vr1Mv0CxgcyOfwA10W+fjxUAtCEz2h6D
N0AHo5RL34V3ovQgFKvj135EJGZ4MAQ/zHzBhOSVR++cnHsdgmLNzA043IKeKQw+YuowO7YhSnbU
7gyZiIQkF00+CamT1Q5AqJA/x+Mnns1sbDS2w4t65hxpm3aOqbDxVU4GHj3gihgKnNuk1Jc/xIU2
RjJa2ZTjUsv/yIH2CBl0ulnVfMf82jEP6jXBZZYWINrlygQKnAB+mkTlelHgvG+70n9OlXq6Y0Wu
qbH3cXkdYndz1uqCuS13w6cTQQ+WSMcmfz6Z87XdGfxyMjmAdYlIk9+80TVoGW/63wMCX/k3W0vm
n9KDrqkVjTebPKprrElRH/EJCxa2cRFlgEYQC7W3sIznQNFiaW1mD709fLJNcgJwN6yskKmn9pH1
jA8xb5Tb5nynHxVxNCPmM63PAibv9zDxbwVv6EQTKRyaWnydzJRgAzPuLYRu9Xoz6zvrwWWZ8Sjy
rb3nF9AgGhKs/xJYsK1WHzieRa/FqOTpCjHI54oLGHFDusHMI/uD20LNkZeySvXPfGgtZxdiK8U2
bfUAIshYdWpKSNy56mLlbakhaeD9M95GK5b6H/PeVbZ7AYpMXFyVBKahVT4NTyTDRIqnk9cwGRm5
hbGpEEl8I3oKQq6EvuhU8iDLsJeaN00LDwqy06g+GL1A5a0Ui9UGNwil3oVLxZSJTngt+awqj4uA
vtgL6i7IjwaxB/n78xcxWajuirF5G9LBiNqApbLXlTFM76nuImxelN0oT5OiVJuafez2OvQt2lFu
Ta8hLom1M0/VJ6cpLjiEXZE0auqA5YcUmXrcQVL1hJyla1ObxdeDW421Fs0k/GqnUGMDMcwvSn39
O9hVCx1B8D0ZL01rKrg667OLkxozUfRmLftIbBcqgqqv9eFTdemQY6tWtasfU7DTjngxBqI/2s/n
p8G3nWHg7lRe1EvSLcR2RSeYe+J2TeSNbNkiQp+x77SH/fZvESAKuKinFTSdG9+3imB6VT2+u+ZY
J8oX8MJB1rz3dcN6nNnViu4OnmdO1QiHrA2d+Iv8ZVutY5OmAJWWWnuy7kbNNhCyTqELzrjmwaab
ygRc/RQofT4EoLJ2w8nskTr+OQBNT744uryAx0doedfpUC2Kta3HCCoTaXN5yL3t4ZpMKY3ffiUM
EUQAP9VPy/H7zZsAxN3DvH9QoYC04E+64vzDePG+U0nZmmVy+bZ1PDlq4CaHIrYhet4SdcW8m337
xORjKdh6brmw+PEnoQzRo7jeb4DEw7tALEN677WcwKPWJBfv3lMmLw7cSLVO8+OX8OB9aF8T93bI
TMkoRc756hitiYBgkrj2IP2dyV6hlBd70UczEPGTd6+18PzACY4wi99cxv+GdftA/JsR6GBg766x
v7q79RcX9BTO6xm9uKJRqMvX4/zc4WCXZC7U7yzC6wRxnzMOIg8wLNs2LkntqCmj+pakz0MPBLMi
CXr0hGEVxE5AAw7ZtJoICtxqQ7chhLbEZz1XPUAmHgYSpUL7mch0o7w8dqCi2/hg0SfjEqLmD4ad
qpwlJTaYPVWlRbEoGv4oL7HDeSGJF8XI6x5fit8dJtQNix621p2W6C20nQ6ZOFMEcD0GZxAcC6cg
2MWAgJWiNx7cBq7d0XrrxktETjqkvp4yp35OxneprVJJp4UWtFUr3rOi/13EF7aIay6G8J1CRX8+
NMep5CPNvbqdxexBB1mES26Yr/Bz5Z7ObVftxbmvYPByuYp9jQSB7SU3dkJbcfdWiF3MCn9DNUz6
P7xaG6FSsfRDz2aE0Qm5830KdXaJVhJuvWt0+McT1vNmClO/KVGm1efIKGK4vcNxOtrOQGrJTGEz
meK4VA+I7cXM/ujGflgXog63IP4TlXgyQMaSuDUqssk4BUwLSxAqmXhrDwrRNo66Dl4sBWAUtl3Q
ndzeNvdkqhN+Nfzg6Jp3N/erGdqxSWw9zAe3+juALJhBBU5E/smrFfcEBRexEdLei2RXCb23zV/g
yyhQl8+c6i6IYFIYzkoXFlmwG6IZVuS4TqcTvwWz5S3QesKkLE4e7ZSrGEpZ6+37+ZJ/7g0LaixP
pvB4YUQHkTVWw8uG62E/icw2fLERsiAk9Crgmjcb5eBXdy5Ikf5e/Tjl5wwxOzW7ueqgGP+dZKUG
ww/Qt+xNpbNNGvZotVZhQEvABIcNEinyFgNEs4uEPaIzlalvTW0a64DT/LHpy2ftv11a5nssVJHy
kzFyZW9YO32O+GsRO4OzPrZB/xe+bK+PNfKHLrvYBhYO1p7Svx9rrlYvITV974H2b5yL/7Lfrox9
O/Ux89l5GQZZXZ+tBV8xVwKEpdBn6YeBERULuHKwxI169UWK8bZUpUTPFx88N3wwIJNhLJ4jIMk+
Aby5KKn0c2E6yZ6KR0162K4J8ayRWlv4l/Bb7L0d3Io3lgqCI2vbzR0+l9Bj1BZuHXQRQrTyZzBh
wsOOJ2qM7HH1mHhNJsNhGbFgJA5wQh3jYF+JDuSpIDJUsNQ9f/8irE/K6Pw2SDQyJYke8VIV2VZz
Qs3Jq52dk1B/TAVKD8/5CUUg65fcMK5kv8cMmx6Vz1mnzQWwUegpMb3QetrDAebbLDfgY2BWCQ/e
xTaD3kECJVigpANXqbXDtR3Yue2NF2RcAnyUuEkfkdg5Sjy20o1SFmNoi2ZyPDVCkbgp78mSbUBp
/Oqmfx7ligwwCOuhfs+tbQs4PL50ZGaq0omQIC9ZN8qLyakWwHA22VlkP36VCytSVhtX/tIULsdO
E/xR5/0qiuQNu+X3WCv1tf09IYfHyIYZ9qWKbGQxahsSyjS4Jcp7Jg+5ly7OxgkcVfX4nSeYLQHM
p4moBFb14Z1ufV9AvI4jfLEdw4oEg2cTAYei8bgZbLoJoT6jM+63GuZXNjon1HMhaixI+WCjWs/D
MBBSgvtsPW4rDNWRx897HVoCqkE1cHdJoTHLXNnrRpQSsjWnBhAaWU/POkEQRsygo9RnK6Enqy3Y
wqBGRH9CR4WXzMApABIP1HuMYGcnQ1bKTZ7WN9qWlvTjcDPFqMtUrMHYrKY1dHJGQbTcIX/WSTiY
Xh9wtE0GeCLUiHRJVPZYiKLrBTYrS2uvrUZ/obfWaItbeJH95tZiIYI603VwbP6l5PZJEZr95aLU
3/zsf0BzMdmBUN10jq1iLTjHI1vHN/EFvsG/DKyKw6hby5Zrt0JP4fKiElyn0ukND8M63z5xyEPk
6gbljBz4bEb1ImMlTNfRTKDpCm7CT4JqgTHkxN1aLg7vbU+UCdeMcnRaRRpvMUA5ITX+qaIirTRD
dB3Toyd6TBW1bxqrJ1WREc5On/Y0pOlpOHmiYwmBid8iQeUeUJ5D8yYdVrgaP82ekCYBFVrKam6J
MhsKye9ogG69nC04XIFWBek+R9xuYah0UuHg/jqI0kyeHchQdCBeJeE2Vuo8YrRpnb7eVwFH6fgD
fNPnXy9j2r5aWN4nXZPDN8hALnlNz4dbAgqWA5RoA7cGshaK7xkhyxT//O/jQwMXz9JKFjH4UhZI
fSBTBWjTXUE1UJKYiT+YNW+DeGrNCLXnlG5VAOou6iYOkzwy+2yh/yeo2YGhCxbJmeOiG6aDRnuF
/U6CiV1LpRBY0LKyfUXouRX0x7t9EmqDlsKoMdS0Fd3+SZDs9FoH0rz1mx65yijr3HibB4fBZj55
xtME3S1FXID3IWrM+ilwNnmlXWO9BPBIdTh2tP4Q53Jn4bSC7b6Hip2bPo8+cBOwcEILhPUVdOl0
Y1SJTxYdyrw1UK0OUMp7LfAOHkI8a2ddVu96ly5o05UPUUDwJcnzTmvWJV784sL4WrUMwkmUctHe
H3nJ3PaHJypriI/gY0a8FbAlPLuCiQIgh++UBiQcN5k3NPqfhU9xZ4dAimubksPaX3GqtD4q6kVr
i2G6ivdgIXTNIKWNyf+r91QjivXRmzJV6g4rCaFiHHGci0LMAJTSCsJx4F9dDtid6lu5OK33ptFm
EPtujhMAwwGIgaFKXnSCRF5S3Qj1oyqCgrS+FnEQiwO4/gT7u33ZegQ5oDcnp6Fm17R/z3OnMzeb
aZZposlUmbllP8u7KxmHpGW4N2CPbsDed/SY/mYH4rvCC5D8RCc4LdN6w30stGk3nbUGJr+fK88Q
HOL+slcJsofvOzeRUr6stFMkQDVt2H8hth4lUT/9iC3U0Op4UQYarEK0BvwtNXDFeKL01/SwoJMu
BtM9LgCb+AO3baUIpAxPgE4jCndxqSC59KwpieCImXnB6jc9Ed4ZRrRA14AGTrBD16PeiA3uEpei
fgxSYwBoGCJxn5PJvxr4RP5odaF70dwnm1TtP+MI08KvEe76Qe08XIeo+8jmKXtSazOpJAkI7xiH
nPldpJ0kSC/zupDNRk3rPSb4wqq8lvL8YAw41WulIdDP6SDRhcMltYrRVMTzKPcit0RNonL/Oq18
GY2a9F+btdK49X6DzIimdRQpBCBUQXazSwm7qI4Cnu+TPSfvR6uR6DvImobBoEUEVDZm1sEgcATm
sj/clDCPuwon05PXzPSo1cQtKljWdt2sdq5QuEL1Q+nzZuaUiuYkJDvloRTUr4U4nvdHXS7mudwa
HT90nc0eYT9QHym2lGD2JWrmbrY8l9chfB/ilTRipwheL6WqFAyLqkiEU4CjPxjo8G6TJtqXSVW3
rPcDmHE1P1jXJtPu5R/GJJAeUsszBfIBD4x3Wm0LjG2qfiZHJrPnXKrguaMvqx7p58aYGwnhP/Tg
AWuoRIclJ6wq3+N/OTqVglfu0hlm48Lb2UhrgHG0bS4FRGhG0MsgdqzvTIgZKrLwWqhifwHChklT
OrctUG1ZiWm4NNwciJFEqK5MnjHDfhL1Ku4ZzMalHjHPg07Jx2Vd1jF0Fmf/sfbsUCX0P4HJR7y4
i8RERc2jBa+AfA7mOGLQjoqtT626GVl7eIqi6dJeMUPw1KGo0Tyv/qORcFf3pi1PK9tRFnlZ5Nlr
wyh5ZTCAV9spTBEcsDK0nAMK1V4zT6YlqnmdZ3LsaUk3U1Lq2FobAkFb46UHLDcq6cRZtlNTMwa3
v/II4da/NZOLxZokb5T6u4CQKFi/Tco5818Ijz1uTLqPYXl1XKxOnsqPBK0f1g90aXOly3Yil8xw
4q7PhjJQO3nHQzp2HEUllk5GeO6CKSdJ0J3vWPTK/h71xQKeMJ9uJQam829xAO7jbCm3DhQ1/PMj
xMsBcFH9dqAo6+562FRTekpiN5AY203EWE8n4pr/rSoPaF0F48r0qX6aJPu8HR6i6M2nvje9DTyx
izW1OK9g0sXpdulfQ7QngcfrK3gNuNfEc11+10OIpWNgOTmcKms74KjsU1NWHX70E/3ZXUDf4Ud3
RI56wDGYyJ69Y5VJ8GiPphy2o88vtsLGiDcdMUPvEpiCd0q593342naDIFHMomBZTE3uA1UgY2c0
vg1LbSzKiX4+eRflpTjUM3Vc3lAzZKMltnUTPNXmpjXndI2KRpFh8WBwEnJ2FNFGE5JrY5lqb7Ou
q7OZDStOMhyGxXKdUiHkkRhM7+zbSCyxsXvn/LLqNBG0G5qF91ZPvZpp6L9LMDp4al9/RtwKRJlo
WfzC3iB6q+ob9ny+Ki2yHs0npHfpTdxnAOMXpUg7mUULlHuN84cxNgh+5np3qImfxRqEMljiUXJn
GgvxIsQKsZNomlmVOji4i9Bh1vHbzF10zA0Ho0Hd9mNAsDFLSIpeMz5ur2QbDxvuNDkQEhLjlesj
S9XefAqBourx0ZJAzTlMNcRioBLCztsbGCvhFy70Psvid+JleW1yiarRaTSg0n8BqQ39Ch0D3B49
QVDYuuHcIbKd+eXo8eD0A5OduZOUmgZjNwKRJ7Vd83m7Dk14/YfG/fldDCLh1ai6vdpOlY2ucZzR
jW91h4rXeIHY32xDI2j2ZR25PXpON9yubt4yjVfgKGBzmgCwoN4OIJfihNIs4v8PJu0WKrS5m3p3
La+KGdMQB2XISDAJsXOfvLAY5I/03DRya/iIqp+/X0CfOVRjza8q4IUA3U4Xp7i3lTP7eMYwEg6B
GZD7URDtvelf6wuCwyz73WpR8BE2MkjipWLdNfItjSg2RfPwEIv7nAYNzBtzOKRdSib0E21inV5v
DeBpq8cADLrcUOxR06HVRPvrZ4ewj7PYx/SUT1obxAL7w8dyODzO9VJmg9yZuHqJRBg8DD8ekKbc
jQSngVlkNfCMER81y+ZSWGXRMlQEI0DVEMoZmAsJm3QA4TNdAUKn9PSQDfTiRz0ZK41BTn7ebRJb
cXHFR/2EpsiItrcq7EVnhuFmG3ngSQrAaE/8QnaxrOgqKGAcEtNXY8H+zv346n5owED3auDUupPA
Zh/aZKtLTVqXpK8I6R683ZZz3qyDjXKqS77PHqwXsASRMJsX8OMKZU5fMZuFNOL9Vm4xCtpuG+x5
+FcVU5hQItMRUaFMJ8TPuSm1luPwH1FcskTWHqAwK+JMVPjQIX9uw0JmnGefJMtOL4z+7EzT0N2b
xbcHUy1nGXvL8byjjXuB0stm35OCDsGA5VJhq06im3/0laY7/SH+KvZD0CQGADPHR5qlqYOApUgC
bbdLV11qGef7bnsC0nNMZWH0IJnpqpYpYDSwGQJDhA6HT6Gz+QFDD41Ciiecx3dhjKxcZ3wA0B5D
6u+G0HeQMDzJm6dq38ODBFfH4uhbJFX+euZZDhVlHXAM3oRuianf4/EUdIpkNsGCW8yGNluuFvb5
7RStnpVkWgtiOt5E1FrIoNwHRZ/S87Iw84xZMlnGEtxIr2ISls7JIBKkanvb20qdyriB0Uc+ld/O
95icHteozO9NUujQUBC49VGhBdOAYoKprzu8kha3cHzrWmmgnAyu9hzb02JHvVNfAIdr3sYRhbdD
CGg9zZPiqsPTSpJzoWRpwcBeySal0+AYbPb99m58PxLArvMpXfOxxfx1DlcB4JR7V495FO8D8Nmp
iGSqFKvoImJLLtH0LxrQJdFVRpxC/vnuwqwWP4jpu5KI37/LnqBvCzgX3WTMnt72rkxv7zxiWSTg
TRTgBy5r87FfgbAtWJOImN5WV++Rzv5HC6CxoDVqshoznEN0XC6jtZl7M0ZBfbGhOI5RQkZ+P+ML
tjsU1JzcZVO+aEHySetJpOuog3TB0BldVW7WXbjfvK7dDulaNb2tb0bRrO2un/K+GEPwGSWjYAMC
Zsz7VQgziBl7bvKayvWo3+YTNzB39N91jBvmUbf7fsHMva1hIKiDddnqfI//LX03UuRA8pH55jzu
jdZgmHrBSf9NR8gU3Tq7YAof303eDsTTjkdMLMv2OVIMt3kRDxGmT0O+AyltbzxLFv25sraCGMyo
v2FNJ94UhK7+a/P7xzRdOKvpmfIv/wthtXETHJpTEu4xAOGyYSaunFiKuv3+pHSyfsFv3XHL9FcH
INuMrXAulMaDqerN/mGW93YlrF8vZp1IdEAadJDVZqQ2Pjgwe5YG/qH54LKZzW5ysFBw3GHK4EnF
eC0xhdj4+R+7UK8IBbW+ba5g06yiBJ11J6p37gMGqF/R83S80GEgvPQwGT6FqFVJ9KCpai7ABfiG
DJ5AdaA9vOxNkjbSf3sGxGN50gzZMKlCIvKZ8z8T0BhXvHAHSFRaqLaL5ZDlX0SbSENN2SZPfvWI
D0pforKj70PlKHagMZJeWH7qs+lDQCqjeG5GCycXYzlBwGvDZz1JcQX2zYulvsxg4CILTBosEhpA
X5LhUoZPkHgh8gTLoPASuapnoLK1kz8x0Mx17SjnbMIExIuaY9S0FhGY+5txqkjzmxG1irSQrKhq
dlZh/qGxiwyuoizRyBl2LVlsODTqZjaOlg41uWt1G/0SWkSjGP/lTNFi6dzYnRam4j01eiGom1YB
j6KHZpMYaOMePtVKN6HV5m4EFP7lIhISLSDsIsMO6rs37OHE+NQUyI0EGx/oz1b9OFPAL3zcpwxj
DzxcTTeM+lV66yMzQbxeZzyFivXImkuYf+KaybwQOazbnO2TQx0Ri3reiAwxcbo8p4tL1+EvjMwy
eDYlPsQBoYi2Id4mVYXXdI/VzcVUTJ8YYllQa4cYJVsL07ZCG9qSrdApDWm6+f+M+mISEu6hhhlF
w+aGlEtHFyT2qEpOPSDFObG+WIQHVJINyIcDgg1/rGAJBTP3VjNnz6q2a/M/fY/Mb8qN6021Yqqp
oqCKnVX6iNd845h/eiLe8CKK0/dro7o8kWwUGmLpcacFcF0nolU2L47+w+ijoyJa+bbfaj82D2Ev
Le1QmbcEhgAtMDpZb85PIOHwB5qEGgxxy8ke0jMxRKVchIC6IAYDImOezQxnqe4P7oiM4tLuYIAO
5h3CX5/4Zc2buWd/LCG2Se3Fu5ndMQkIEwEZoLA8/wcApl8sBpxDLx3WikKVpgYXKuncLrsmdeC0
9JAnANJCZi/QwT+2LvHpC6k+4sEpGZtaF5r2h2Tgqwpesw1jqAZM4sEXECgCdCTLOriZjGvDgLJq
T+CIwb3wIBRVOsenI+97lLyuem7EmdV81oFWaWH9F0Bxc8bLiXWPucpTSmOSLyehJedj4LgqBb6Y
c49M712kX4mbkGWzFntZPP5N0qZoNlB3d2ZVUDID/oU961Prvf83ZhCui5HjK0y8fEXJOw65+Mat
o/WG/fXXerq3ueKgMt6Nxowrp/Kn8j8/3a4CLTxzdyh4om3HWTpdElcJzM8DLi8a772msWcFkQpZ
U0xfc6KtdhJTRPUXcnKo+87ZwVQDczOTL3U3b0hSYM4xlJoVK+gmPMH3fflMnECH59NbIjymZ3bS
R1bm4iHUpyzwG/UPhmDLfgNzBXk8U4LonW5/0l1WqfuWNO7kww2hmwPDYvMaFqT60JvHxaAueT7b
JcNBRuh0lhYGPzDIdXg9d0QSqIgs8ramON/3MgkEVm3EUvBxy9m+TzqQzwQgt2oeaBViVRSm1vSN
hLEOK3IHuKBjJVvLBcFcv7dTJOpsDKr3XZ1yRY0k4wn1BfA3PtCQv1qZdk9G4K8gcPY7g7Fm/OZP
/lkk/ccUxnraEhatTjZ8Z3e6RYUVXlUG1GGcSslGXdCYxSmla8klf0ydkC2ntIA5eZA4xIRhULiK
CTPNa1Q+cyP9zuBSQggbOwjJnAN6sFEiLOFKLaMqjvr5jrzCRIzJxnZe6wzfaCW59xfEv4fTgQVb
HyyxvLQbMBVxUJVXoO5BdxDvzJyr5QsoFZiYc2cPldKihEhfXwclChDeygoHyhxP+xeNoh6OK1wI
lXKkiiHUVqxeuNXIHMSl6LtS/5qeOqOAuFPue3f7otIZKtyQknin0f9LBn5WtS51f4nUwIT3RM2D
lpHIYy3tTFFvZw3kiAbyIZWlvx0WFS2hF7NTVQQKx4ad9Xo1kgXbU5+XpMezqnS0dm+kZG52XcsK
C6W7QYgqfoJZ1w3mYES0M91k2XdOu7uijvyzE3Y2L2SX5MysSUXYmMz+ujyjYw8HY7odBUVqERT/
awMYaPZAEKyr4arSf2k/+oi01zgZFf6Fl0nQFdp0QY/S74ivfIjRp1x5ZTSjeq8e8QFaSjJ5D394
EToKRjqH7VM2CUtHIiB1m+oye03+3V8I34hIjhxSmW2e6mkaY4vBjnK/7/gGX/cpTum34oP+LhBE
NvcdiTTmLbmPeevKySYYOTnyqTuwDmDDhJxZj/+eeDvMIkco0Z2TL2qX7/cEAU9C3cD4bDASUFY3
y5IWr7Y5FUUmFnffaNi7TLVj8fgVmJBOtnSbDuhzaxz0aBhdg14/3Q6fsP+b+tcYgy6CRpROU16a
3A1WqoFfAG50l0XHqTiLpu9nVJkF8M3oXOURVVfvQtHNv8wL+8GMFqpuOi2gJmrrQbRzzWztWbgE
kr+V4Rq8vHCEqKPvsukkkbaoRyenXIEj1iB7tspB98Rb5ImVri/4ossBkym/OX9V4Efw8HuLD5Z0
tXFVzoEhPp9NqbbT99LacbZzBMTSOPNwcxpmdzSDDIC+Wo2Q7ZtxBQ2QTr4uQxMYkpzyOWYKoX2s
I1rwFWC9JRu7czQg3MMEJprWq8UtRnqzUZcvC072RSJRblWoPCCdZLKWRMG+mvK7TKg9IE4F8tyH
BlTVv1XMgsas/XgcxhH/pQnqxC8haGQVflAcw+/KyXlG22r+FQhjITqRYz1JCgJjUwHONuJMuuOX
c6HNlJ0ht1NmqNhOfZwqMKtk/0Ut3GMI4e8dv1dL6Y+RY8T0h2Mb/j6TAqycHKOCWOQt1KYy5eec
F9ogvrdemyx6sTTV6pRKeMtEHUR33/forc0u8drTkRkvDYgdsHGeGdkk6ZoBUQjcyGKUYwmEEGEp
wNXjYGtO2Y9f2ejM/guQPHy0n8SsU4Ly6y0hS/r4AmVOh8p7p1YdM+YFtONbVNvLP5pW+wt9HAH+
gEluhem3KqfjpP3qb9DQtbdZ7Pjiy2hyDFYvAu9DfdCDK+5R0ukGKOu+fgyYcjMQ/uIE++/ccIIO
sHETyZZFX9mJ7AmCErS9QBjTNjDOQ+eUTmxzieFcVotUZSPkBhAfRrCtGSizs4gcWcXwnNX8kNUi
+NY3s//nzBC1D6bGFgVRynhMySi9/Px1NMLmp3F15uwG7fQRoSonSPlZY9Yt3hWaQFWywYzOtEVG
17xjfyfLj+jiQpGXhhKs8c5hL9KEs3Py0gG53jIZzbi4CWNuRXsWljb7ImwUdjVYVNpSbpw9PhOd
MOcGhXstjTdsK2pzq39EJUIqoT8XOkRrsjyuZ9nkiS6ANY747PU8Gh3ril/XB/DXfs1W79Ejbz5j
5kbhrwTTnwqJ8TJ972tBXacEJky6qgYNCvbqkkrQTVvMh3ERY2k8lGFTOhGjICe1ESl07FQnNp0/
p7aGfuzS6m15Dt/tS9f7C1RMpOSi2fuj4DEm7vaVVJPg7BzwTGq+SsQ83vEoMs0bqpu3AH6IwS2i
GJ7UyyOHDfVJKRMudcZt6fg1eaobYu9mu9CY0P/RgmX2EoPoqIdYr3i2XPbF+qzaUuiCCCOZri/4
+Bqh3XH/tJg2kZGgXx6gIv4Ujb02opiUEJSUUG8Bk22RVuS/DqrCnIX63U59d5fl/6sdEFfnrca7
dpN9RkU3N2xRBhpElqP5bbJL3ANixWn2pUoS9fWC1R6SHavp2dEOabrhs+hZZR7oWKVX2ILym/Xi
6C9KBtFu+ihshjM8vqUN08mvX8rKjJzTPWnFJe1Yr542EAT6mrsF8EPZt8J+PTu0TXcQyVZg1Cvj
ivpIFwdzE6pE2Km2AtclFpSmv/bymd4sj/j8spYTSsbD6nwPqZuChL7SaTNrqeq5BLs+udmxCTDA
645F6YntRjAv0QGhlg5EltMEeV5tIikwMlwcrX/BTIC7084JJRUIBhhh3Cxa15UIA0SsSBRG4SlN
nV5VnrCmFe6oQA6vEaovpumRDglhmPgp/vXthMfG3AEDOH0ATo3/MAdCHnJojSziMMnosriuO4jr
sz+3Y0uPWrZlH/DnwyayPIG76WH8G2jfLMKJ7KX1xWIgoYMGFCXqd0CJYWp8Vv+81mwMpK7JFwU+
kvhi8rJz2PIN5DXv4D4pHC/B1+t2xiZrHvBL2bfHT6u33akM1/3COTOngXvkFyCIr3/sKCU573C3
5AQKunD+oqGBTXVGF1tUyav+Zfvfb/IRTy+H4wEuyiIpopAjOO7o8FbWZj7SSEq2hZaoJjqoWUyR
EHa8gp0xJVboZ8wJv9c3pum/bOjRDjgeGZKxWPwQbdSw+LpsFvt1wHIjUh6iz6yC6rjRSEO4ngqz
w8/BT4x/CBf/jU3o3jx7w79alYtrWKTv58Y/XEjCGwlnN0T+5Mla0Y4jssNrO2WWPt7n9CJJ0Ci5
YwrXHNDx6Ksp7iaCC0MSxqTijtRQwz3IlZ/ejib7voPqRiv8xfJRWVstIf3ndZXNJpcutikiT0pr
j7Au8lt8Cc47xMf17Zd5EAGz1NRLdgpp/qWoYyF+qrMbY49OmBU6oMQGbCSnc0bYAfOxE+4ulpaA
Hz/PWxlzvb2hn+ondyKrT/pCEg4/WKjs+355rO8WSOXqPJG1uulHCuGIUhQNByuqEXln3TTEWOM5
mAZQ3h/8xe48jcDp/ZHn8RXRErBxNekYbsf4VHbfYosq+pYAJJxj3ElPSN8lSQ17yk+MSdVwvl1i
03audFC6rSjYqUECxTnTa/LmKQMufhAVUYivFjffhx2n45tQDJH7BsCiEKsfgQIFDjx+gN7Oo/Mt
mb+KdrNHPz4qtek8s7s1oSG6dhDwFUa/n3P7upOrjl1gnBbcLDmDkRhkJbUvmZWfJb7UMVW3VUmF
1Rx0LCuWOu38fUJceQk7ZGjMU0q8pVJHwE4ivKMdAAAJuDnS1CpoVm13JANxgMcZ1Z62zmm+RymK
ymYFwhh6v+z6760IzuB5xeGvBirgQxUis0cBwek8hGvPRbqbAhmkaVTB1YiuFQ3ZCkOLZEGENU37
97KpVyKP1LjQMivCmBskZDz3T2VvyPng6mrX1fVc/Pq2QrVWryFdbKNd/5ZUootv6yS9KGJo0LjY
RtYiNNv/LkeJkJdBUbvdJHhmqy4xI4sqtdxvd22cnqq7+5okqge6VPgk4d/0TkUCXiL/0qG9d64R
1SaPVxZAW+puIt5CCc89x+TxgAdFsB37inCJ8yOM0NHffgX4pB6g7TvVmHXiweKotH2sJC0uLazI
ukxIKfN1uzm6fN/B91YZsYcnLTQyoqlo4GZJH7H/lBVxGHVEha9v0jr0QSdHuGuOwAmd/0auitqP
Ld8mgJte1MN22bIdsC2mQp+TXzf589V+sx+DlxZexueWW/o4p3E269p7ftoBPh82fwRQP1uYSXAI
2s+DlXI2tcdOV3q1oYqP0kqF2hJ/zoTO3hjMo67w3Rhr43o3XEBI0cJAWoQDpd7ZdXS6eGbR6u6U
YcsKW56fbGe1Wps9l69w81jd+zDedi9Vwa3kpnxl93II6Q02VNe9ySOsgHZim0Da1KXz6FesGvho
mMX/xkUuzlCrIK3DcSyx4xgLA187jPv9zGarfopLHp3XU01BLWtZY+JcJh9EXNXn3cah1o8CAd8O
yIYhZri1dKkwuXc20lJ41j//zRzB8bqKg7fZ8EIIN4wYgN8GuD8PMMQ6GrYUG/MDjgbxFut17FSI
Kpj5TAuPyycSQ4MmNMBIuOfTStrn0fvySJs44YrlkCuXgt4X9OB+mB22QAxKa0WctQYFsgbhBz1K
JI3wkjCMp1ur/6jGCWOw73De7UUaVlwYNO2Ov19tmsLKqoLXVyaGq9MmCQ9waFwN1Lm8TpwX30Hn
CZx80TQhMKV83T9kpnu2NypdAMzmQewYPfWhAd9Eh+eXpVK5Kxr4qWGgQYHSnD+1FWIZHkn+3J/I
7zYG3Ghjj5qz0zJamSY87NmyszD8pDjGNFa/offVwDHBFs4garJcEoNcsmDesYeA/0dIN1USg6c/
K3zNN6ghcuyUx12eZTWFKgltk6/BI3xHMJWGwPTr+NQmb2xACfRNu8+fKC223vOkRIbKjGg8c7rM
LhStXJbN4b3l7R1fp1qDrnrPaRaHqunLmyu9oKlDT7RwF9BqHEGf6Zhk9Kg9yKI3RlWKWu2abphv
HJgpZjakNfo+BWrzYVhbgM2awqv8wyuHBwD5VXhgADElHtSmZ+5Ik3VlmsdITi25z+S0zzWqfbWv
nxbhuiiHV9+ndO94dFRe/wheVmoJq+M2P1vo9olpDTrwOz4iKwXXv9eHb+AYLOMGL4/dqVE5hlG3
tn4tBScmIQrvq7B+vwpPsQCAl/+SqRXkLytNqPk1iLVEUT6oiV7NCqpva6Kt5ojHUJFXdrhdw/vx
awSHM6a73FXlGUP6rhal4kSy1nrICkZDiNYepikb2Yn5WQcy/c0ZdB+XSX4eFvGGkSrmHdNRpGaS
jSv4+DoDki36uMAjeKm6Vwk8k6XqmHZpYMWVuBENwBeJtsC1E7yjgv2eQoc0I9OUUqqlYOCC8Jk+
8J7w9SPdOgntOUo8y1BnuHngdYmL/ZY91Tw+/COMMMdz+HOBSTNdJAf8JZ2+9M4ZZG9dcGoRnP/S
mnw+mNrcLyXZZWmqmtmbFxVjDGJr8f47hqEH8/xcndvqyzJEWNatYcmGLvFjF8/IxZ8snSLmQwR+
a/djfAsMbIfw/4DOm28oVvo9wkp7Rc3uP4VnC7KzJGROr+scElWn1GUMIpG+nmvZcwiV0UryZgJ+
9hL0hjdMZkokUu/i01x0/vY4RZ2ynYQx9UFcy7fbQStYB5iU7wOuiYR9FMaxN8YtZTnH9tJY2DJa
hlrsrdFbKI1Y6Zp6rwiHNkwVT0tk28PuT2XxmFcNpR29XFnMGSurTXsb9y+YvrLJumxS+HRfpnJ0
UuARYMZEKBwb3SYzZuhBHXqxcA/rJ6nqhF7tC9aSME5/MCzKLZMqMv6L5ekzxMaqQ/7n8ZECYvAN
xlaIRwF3bFo9B+smaEwBIaPcdrFPpnFTmuV+9+YWazhGIZG/pYgpa12FBjtiH9CNz9sydW3rnc9H
Ydh+y7iRy7+71FZnPvSxZY70ABUoNLketUicHmE0NLyT1H//SqTzAs974rUJt4S0RwQtUanAyKB6
+8uQSz9eMMd3keltGy/+yBv0QVsrXhWGOpcJJXBJ0Qzaas38PMDSqUhjJgtUf4VWoOqpWILkEdUf
tsEhucQ2+i/QhlQmqiO/6+9UkgLcYRqr8FxY/t/cGpHmWLXgJmpbIku6JP78NAInCQb2JxfkHnDh
ECFAft/VnXoRwqAHjnP6m7qHWiiVnZZ631PJB4cnJ5I3Pc3d+yzcuE3/0lmby7Xu7aCqfYOKS2Wb
NgdjXI1Vni1Q6DADY+xII6ESpMnT8fsuUpqaEWB9cUeFiuORsVXDNmUpc7rjJ9XoqcxxjnXkl1f7
33btG6/2XZizlzEEOQgau6mRieVzkoAtWUKDVGDQaC+/incZy1BNqeyuhf5W9eE70CeAPoeWcY6p
C3EkbhovwxzdzJ0WvuaacS80GfsoWjHYxxniugT/MDtbOGCA/1fh8/F9wbhgICsfh4Dds0jM+Y6p
rxECxSelqMu5ylV0cbloynZL4DnkPxHHEsFIlNiDOAIueWerbiLaPtQZJtshRMAHB8wiKiwxQ1+S
+c6BO1ErJhHnVX63lydoUFlwn/QK0sgOZbN3mMNVvYNfvKp8R5xpVDlfEQqYf8wP2xatCAICRIAG
vvvhzAUnzikh4jqfPF9LhQVQKzzxSGzN0pTt8SBqu+HX1kZ2VixR5iaGOzpUAEFL48Ze/i1drq8W
PFSIHx7PD/L6588jJ/wFD1sT4u14/1gEcOM8TP1j6OSeQug3TrPX1bULmz5GbaCMV8MpvFaq44ia
CoG4zu9NR0N9oL4DU7eq1ymEUnAR1Lr5llnCd3GwwNqjaHkh1+GzsqRHWxlQlQuP+peZ5ODYvpHV
/XKoBtF+qFnNAQ5jZBBCk9E+Cb7U7alaHGUUj7gTLYpzJGmIBK53yB8FBGb1Nb47Dd5J4pYi8cSl
hsw0z+DqDmlJcMiZlE1L4u6+0XKQhArqqHMghuj2ovIx7IgqXXVDgKsd+xPMdmleYngmEWboNiuN
zXu+oHtq3oqEEisYIGJ61mzFEaOsnhfKkTIcYwxqWYa1RbbL/t0FC7lJUFkv4PFJ5fYpzC+ozpP8
RrQEpUWPyIrIzA2eT++joDGs4/+ek3IS/atie3iEUrwsaNHASedS8nou1ADuRlK1vQTd9zUQF/i2
2xkNdTjzS4Mc91qMIrKeaEZWKI62uTcCn2573GuOEgWpnZ9ift0DZCfyjHibA0jk26K8PWXgiRUf
CQNXnVQ6HcYbnKxp1rLUokqMMlZEWr81nEg5byQdr339sqo7n5awZO5JnlxmzmL8clc/xx2Sa9qA
+xTUjCf0fcWKMo0s7Bk7j18wLTtwbfqa0MR9wyWXrNNRL12T810sCha4iwYEnPcH7kByaYyj0fyG
Ib82zCSWwNqEnVqHk+z1dHMzSvkkBcJuA9O1JZvq7atrDF1zKJeDjtALyMN1Vtya7nj23VKoQoPa
6HJPwp9EAQFDOvHtw8U8VngmMHBC6DWVuwo2mRmJuDgQAMiP84abW1AUas/72qczX25fT+oWe/Ne
7aS67jNcKigm1beqZENt3cmDmSw5Qq0Hw0+3qtLXAm3XbsyeASkFOsq6wQMVxIliGWk/jEQ22Ipc
yL8mPWIuFQeNpbdkC1JKZ83bsxuO6Ci3+/a08ED1j3p9JU82u/KiUsMKQ5CxMncRLsL1Nj04tt/Z
5Vcev1jyHv2liCfzfU/euWHrUVqQFxWJYxGCr8bXoz+nrhhk43gIrXxltFIKFglca/E7By1T6JqQ
mTXt0VVTHxmFV5QQj7r2WckC7LFrPtnIBM+fxA0MB7IFEh0GhbpiMkH0ZDFqpqb+1OzipPZSXt3c
4mUMwtYMRNN+BfVz2dFCNJrwCdKVUgcVrpIxVpw7LODGpe/z3m1e87XPvvbyCN1+rBUtRDYNf41e
1yrHSE70OHiFFXQJo3F5PFdC7WQQbLggQPJMRxW+4/nI3TeuwYGC7S19oHX7NRIr7j5aniK+GzkU
nFud1JjUfEWtB0IteVx9SxyWQZxhN+X11hwxZCJBPyloR+r7Veyn5SAOHVkHOB06qZqg83g90FIa
SWMRGD2IdDE9c0WTUZ0tkGT+h1ZUapWSsot+FQtoT1437Y4OwHEFrHxE3BMMiI70RCHe1ofrRP6x
fCX05MQADgh+lgbmKkG4PccF2QQ8CtzbJNIVlbP02WDlrLeJdyF12qyWCG/lIW2ewH25R7WhzAb8
ehHKQXcV0LyF6agPRNtMQ/J2jXE+greK7DvCNxVMc2iDVSkR/wp1Cmdoh7pofzMsr6QI5UHiwQdg
DY9VKyuVUWH218fwcL2mDtOdh78roj77BoZ/99hlQgTglPSqDhRQuM6QBGps2MuB4NkZ96L/9ETE
1nrmMJwwEttRaGPNG04vNYaIi8SjpYrxUuEUme1KyZWgP9UmlYqnuvMshuDNfG4UIR0zVBXEaDPs
D774EH6vJE6PQoGznWwv3Ic9hH9BTHay8C7Hq6TcuDTNWd5qUNv2gmnNe6idHIlychn5n8emWM1q
RYt+WdiGJdY4uuixrUCpn+YMNVEciQPpkUYqY8M3Jy3D9eQqK8X4LJzAqPQmRyG4qLiEK7e9T4Ac
GyExAea+8V5wLdK2TeKx37oL+QwCqoism6/UfD4wBVTmbiBo1t7eWBTDWTGJCvzRHqwnwdZQLZaR
5u39twIkX+LWy47353z+Tv5bt62sRivKFyD3Wkngo046TxBE4vlc4Vshj5frv537ahkmeJtlDFCE
douWQX6loJIzYJ4CQaRK+794zRjquSWFIrsZt8PM3i4myO3BwKZ0oieex9GYhBt9HtiRmesQTSBQ
/PNij5iYqGd89Xq2uI9Qg75sRVGVzsEHFfU8iA4NS3Ymm8VntE2pIC9+b5i4oVNBr6aVKv31Yg+Y
gTS1Qhgv6YdGcIkYubXHWHQjk3LSVlhh8nK8afjuOiaEzXswTduhdEYLa79MCH8617jmZsvNDU1/
MkYLmDhiaE/hjTxOclkNZq01XsJW0iNjEpsCYWuY7IIRet4mv/WkZAx1xS6kQEQ9DneX9cYaHZGx
QHXzU6823urG0K9r8XEYr0PbCV4YrCHKEFUOI13aeDnCz7vQclRyDvdnElNP0pUOIhoX6XgN2SZs
ZaYcVd0ta5VNiBzNkt82NTdyIS/8qKzZpqj5z4OC84tnkmydEc6ckN72JI8Ym96YYJf2SIqbJXOn
Octfnlq2IJB87uJiGfDHn6WTBz+veBT65L5juY3jmj7A67KsZqhvX0s3/XHD2UaqBMawPULOsBUK
1CjcdBdrsHEuSTIOeA5szW0aG6EcAt7oUQpjQSL6+QgQ9Ufaygy1y6wypU8Rpxha5njmNLpsSHoH
KUHb7aG7s9l9vjmDV0B/cHybKeTTDtf6hJPOs6OziB0ClaJl97slp4uFj3Xi7q+qeBDr4Cb7wF8/
sBkPe/Zlf4ox6rXPOAymjz/fhBHtjoIF5TL++0p08ZchNh8/BuLd89XGxxtgyv0hMZc+V+odSy08
pAfwqM3bPoE9eb+2+zzbTSGleZFlsmPdPCdTPUevtqA1O6ZXG1tPKwlplsKQHRgXGZS/ZSoe9kWe
0GbRxUTrdwRa6ScnzYbo5fKfLXJv48N8yMYnYuOxZZfc8B1LZGOA1Y9GE7+tS85TYcsA4r0pSoBH
+tDKZFCjk8IPPE/ffxKltk4ZPu8hTq9h6Ivvr/ZbsSPwTRrh2Dd3yH0dFS4o5TVavv9r4kqRzEEm
o7rm0eHENb1qNllwK1L8RmeJd/sZ23tBViUI+A7I4oF12aJviWHie/dolTGcUB3uVcpd83D8UgN0
Y4EJiEIXGPSzjW2Fz6vFk4ngF1Ws5JFAsCz0gJ3bmeleR+AJeNZmNjcSGDfStzoK3RMrtt6hm5dB
hj42RmRrSdT8QwwirBn/1Mo59KSjXEYX/vgrGc01/sHpFNC0FQdl8D/pDISxbvEbIoGf9HAKUm6y
ApnjaTyLXOJJ7hACMQNYggWaXuRUK0L2V6RD7+nHsB9h4+81xjPX5clxEFv4yip9HlNMmKoCrZv2
OEMfCUMV0w21uzre7IvGDeWg9SSt71H1pmTplpJXTrlsPGeEWOwmHyaf5Nn7vtAnkP3ARGHn2O8p
vI+rfjZxj+38XnA8bS0ffA7FDCT9THQhSh/kUtsXL1hjXG0foRTeXw9WrckZGVFioteorXEWugaV
KpAapcXmrQ4U560nEQCMIqhb7M4R1/tgczKJFrKMVIDFLXhEHJEYhI3Nw+dqW24VzFmVHuojuFrA
DI2CG/+ru9IcVMDGx7RCKtgWj7ljjs7ko9Ngd3fNT6FDCJ4PCBdDSY9fz0oTKZjKiIgT6uChOM06
v9DjjAIcCS8zo9V2goQrQR8sY8/uxGP8ZxcvXd4KwsDhNcth8EQWWulxcoc2z4NGC8i/V6MyHunx
wtN/Yu8LMNIuTmJi/DyO21bCywT6StPvOsZ5cUPC1LIdXEgpt8nA540ZLtC2Alo+VXAHDZ69Qsug
LKnnpFnYCNUIap5PNdTyJ/7GS7RSwPA3FuwP40Y69MqGdXx1URTzrQhibUa2biX+L0JtKSYrAYu2
CxYXCo+D2xoNF3qslCnlPRC772uXYWO7/BxzZv9LB7/KJjLKGviPgqbyFArViiMv/NrTJj8KXP/k
0RDhdETxxfkE/b8wvoLiEU49mmb0Ao9dLcfgYCAxpZuacSR+dmLj6eQ5IaVhQ4zprsepUEsh4FlQ
CnN91glFVZJg1A71qxwQJIjL4BKQBcfpBJIMFYSPB18nh7uYTtIwFt8I0CvkqMAgBltufGNcB+Tq
En9Y21C8sR9MMZSddZwOsXRk7CwLrYkDw2vuBiYN6L6F9b6iSp5HjDVTXjUJa3ZNFGn6LkBLl7mk
IhHSi55vB4h/I+vGAE0/CxARhhVLYAJpIwUFBAwlL4Q1D+zIwo3L22zHVULX4/CggRBBPc0CivNE
HcAB5SknHY9K0/SrMi0yx0j8ikZLO+2767WBFq8akExjHnb9fHQAzEFhSYU1Y09EdqwEBgoFcBmG
2JWQMPINem92cRJpaLlu+/xLleyMgKcmD1ggtoAxivaS4mEWuFUeYZ8Gs4nDlDl0p6fQnjqLfXeq
g9m/jqksT8B26GtqZfWY2JipKHnjOdc2OFML4u6SNoGW0r3sufH7EtGePGNVox+kF0muRU9rs2Zf
SdmkoAAFXPBBV/SrpG9xfhZPDrSWP5zuxmELfhOeKvhgwqP3EeN+wW4FHaFxNIllsYBcQYWGa8Iw
VN3ClBJfdyjXRdcNcWFfs+15r5UHBeKgi97B2xhlypsjXXBQS1E0mTxgUkXSNw51dS332uOqR8gP
CFE3SRrNwm5HfBc9cDcC4oU++rpYVfs7byXH4L9BRNJ90qS4s4a4qBREJeWDE/1UDbSD0kb5si2y
gOFV8xf142gaX3GU9V5aU/R2/xBxoITYQuQZUFve9MHCg7mHOkhsODehPZ1tP4jkatiuI/mm/ytv
XzAT/p17qixZTlLu+gXRUn8W8sP9aH4PR1AW3f2YZEMzFYX801xPGTpnIQZtpbZrnByhQZDlp6ko
oFG2LrWR1W27yrsVLM6aCPCsDcHyX0++0DaM83iOEyuYyFcHpM98oiX1MkftpHAmlFdfCWfQVqSy
abtgJrjtjVHjZcuVq/hvKXssAbzzMD9iKS5Gw8c+vcJpwMOQ6PhfGHufqw71pt2+oKfs3WHrB0tf
9rs6LwjpM6xGHeePp2+C9uFY/8y80ykTpCQOVseaoCyQkcHm3t7OXMUgKt6DR1gmrUw80q+twOZs
Nsed1h8WpAvUH0E7lB+lOvZNvGakOQs7cxoOGkV0M04319tdIpG9gDR4iaEF6vE3L0UTq5EWenbF
R+F4qm+7GhvLpWhrgvJzoUF9H4DAbgzeuzKOGBlMOul29oBlmOchOdJ91HgUfN2X90MfBmlQTzKj
7zYmWGruNDyp19hqCWg+HtIYyaB86IDhIVMt1gN2oApaSEOidt/S9FrFxpBdocYEf4wxDukuE31O
XecRyRqqPHAD2hUUvZdLsv9jp+7VRmywN2O8zDyU1Mi+1wo7E5BIWjiKU8zL7YMfS+eoWnoGKnju
imR1NYb+jvXPIkowzFm+X/iIOjlwrq5fhyBYyaqhwuRcH9h0anfFBwJs5ks0nIrolKxCGaiAlJO3
JrvLdGVAPIrnTUnmwVRsZZ57ZaYaLJlKPJ+FIwbL2jsJBz6r3qFKd44//OPPTQbi7oDwiYxR5wN4
hRTTVScQJVygTc7PG/b4/0LrPUozXsqHvAbKD8pWTGaKToTFpoiUPI7Gjy/3pkmSIjK9stqvzUjy
Mt6uAZWLAgpm76hwhle0FGe0gTu5XhhdoWuqzWw2qivIQIln3LdDsmFqsVC2CTzsniAF1kCnKF/M
MM9q0JL7zEyy96lr0ojeVALAt2ZRwLfwq4K1R2aRGTf0WZGOhhj/3v4AXSOVsmwRPYi1vOFIPeQK
YCB5TCRnJ9/NgEbSO4CMT4zt5T8PggWgtnDsr2LQCdbLLdHXikEm2CRjQmmMZpkW4f+Fwkmdg8r6
l4TGCCXKpJGa0qGw8y/wVGkuB2I/MkcrQMx2cnZKFexUIzguTL2b/u/yKJLpOIVluIGhleEDL3iH
BC7a/FYx+uDtKmitzAPPWVbUemChasja8DdCO+bFth510LTNeF+WJRJIN2+bsst4uEJmfxPOqat0
0nxSI+vVcTrBzFI2oSoVDptpCVga6pkYiBuBG0UsnnRWxpiUmaIbYJozT6GQCF1oQtud/N5sYegO
PaL2ZEaRiejRymefVYecsHn5swO0Bdc2FuVhL/a5x/5D2mW7I7epsXrs1j8EDShrAju/k6e6k9+O
aTRQ17ry+1+lqtW5LR6mvm3GnSkvpB53hTMzjD5OpB9APc+erVBp89blWqvBKgPA3FncnBsLBTBb
kpfI1/29/ZA4eVolqfkRwMXAPQXA0z763/o/d9h4qJ9HWMIyofeoOVISYLMoIPvWWVzcUaGBVotn
UY12VG/1tS03iafSuwlKrNm9yPwaojU6ZyEEsEJJxLxdpQ31oy/4YInBbBDTZDdJjgNhvk+zaEC5
t0/1sJURyIGxPeeGTZ2To1QQUyjU8GCYYFnWGaMcveDwl9X0Uyi/zkNY1kOz9eSCAomnWfFAHAgF
Z3k0GIk5MRLUF7cxx2tyJgiZ4wB3vuU+JkpyeEaXOIaDeZgoi+HDRD2p4foioozOvxRrmaNYDLMM
a6hM8AC8PMFmNarYIkMupTHLBwklSOViJZYeLY4bjCLOkncULR2BxQFtyP258r98YSWMh9sGXlGq
n+HbjW10F9tp59m2Tqed97Jfgl6ofdYUwmULqHzg1EXrjiNC+thhW9Sq/DA3HAVEiNDC5UGyHNdI
RG23V7WTV5zVGsswqE8GN4WKGxQJ1Zfg6gf3AaI0PyK3J5hGer+0mvyDL8JlOJ7OGWjZPwLPRabC
ccB9Fo+/P8TG8ChcbVD7pbnjp6uijkW+M8fu5rnQcBAPZP94jSH3PwvBGElOI2MeNCjG+bH81TVo
uZwaV9QAfEzeAFHz/+WtwqME3YZDh1KYGxCOeJWmmTi7BcA8hS3LbCAxcfboX0QIqS0RHbeTHElA
wXjxOmENrfvZjey/w3VbtkGNuqDiqIeEms0qcPK4auLkU3KZ28ArMJ7BioEjWtrCuo6DH/aEgwMO
MGnumJQZUwt/qWSDGrTUSO2IgqUJwU1JQUIo/YkRXiXA2j7wM9R1U87p8BVSiO2owztUtSPlfl7L
Dkjm13APUeV8KHGgiUg7B2GVJiX+9tMWCsG5l6gHTFtDv4UOgJtM+Y6PFG8zhDGTemF/Z1aeV3Fb
rKfc5GnMyjO7DX9+/P/o01jUJZAKzZH3jGidmSahI5Lr6Twiblrz5lxGviBMsAqU0eurg5umMh90
MFhFflzFH7QsK1f4k2FfjPldJ0fIhLM/WwrTK2tWaVpIdJjrP6ZsmMwez2pR3C7LY4CQ88auRxh1
DHKSSZ9wzzF6+l887TJpJQcNFaVFBBJuGamtTspfJJFjRjjmtGjuXtKkZOzGXIJo78CyEeDBuIhK
VlrZTJPbzh2GU1FOQ3kXMG7TROLceEwHnbaKHfWsqaz0zGN54d08XYGsttqpusUgzrbTyzkB/nkt
cNDPdEjUwXhve3ESCrXoq6KmJTVPIexy8XM4bVpsHJOTR7CuCrfu49aM0dn36WgtvAyJgTKNeGDB
T9MDcZ3GFkc+xqTmcf5oj3UhbBFDUITwkYiZWFvwNjWuNUVUACtSI902bwPSvJHOGFqZdJhcgQF3
tljiBHzVQC7mpZdspixJiTPARsytRxpoXyMXAH2bk5tYxYGkwMta+8vLRmgkkrcbvYYHegl0pld0
JedwNi32B4kDxRMdyCZ2SnzrB9vnlqU+FQm/29Rj/wJGHjrRXdiLALMiJDFnDPWfISjncxDCBHjS
znSd7pWQjk2LLcRPhxr/yBtukQW7LQtP7REV3e5AjZVlczG9Od2qaQxXkOiCkT9lG3trGBVAsh5y
ak7GhzSuAymdJ/5CAzPMywhdjl26G/VsHMB6MmOAI1Pdfo25ooUToiE3k3SGGlNo2Me1iKj2Dqa/
wg4LvRtKtycZuXaqRZr0q5evS97mLf6HCqabw0DfLX3+qtHr0xEr8seibzbWIXohc6Sm5Yfx8OM0
uLfCbuAwynkc/saWsDaKC3L0enh5za6O9whkjpIEVYngWWhycQDiFWvOU+fHZLUVbZ0Wq8npY1Mt
v+nRQaGUVVUoDPVsGptyhtsp8Dk59ZMMgxzJLIStjRoc2syIgA0vBOg5+ZpWsCIfjXCNMv8eGBWZ
u+IBmHX22D17p0KOYowgE0dR6WmPAUlMaj2DDZEJj6s1MMCYKQp7kHDshT6luhdjIjTEQ+q7eP8p
+VIUrrB0n4Zksk4Ibiz23ulrnWxxRfdNVhIMcXnqdiWwUmxrjo7DfOcLZy8LrsI1Ap0UR3V7iauH
oOG7UQiUsO7548MYyzVRnH4Jt8KY/dR7Hn5XMdV6naof7uykQ0cd2UKNt3nl031pamji62uAlyT0
tRGopiqXCIOUN0rW1UXfipiXSy/xPuJCA38IRev7uuCLNW7VMjtbX14Yfr+Q++CrEgzgso/5gAJ4
/GU6UO1/51fEc/6IF3penbrZv9TVD4nviiqsflhz0ScyjpJcwzdy7EPQB3HN/7vYjnz98JTemcci
uFjfe7DXO2AMA5cQ/cpo17HfYnyG1hv1/+iwfZYh97fo7TdZ5I6MdTymlFHH7E0ULTKOST0BOWPm
lrfepr/UQjd44SCfgr4mNS4Ptr8/XSkRMyuYZeyb69og60tJoYDZtqXuPi2p6NT06uGVD/KoltGi
L2PnWaC3dqdeDFk+hGzeYXxxSnWttcip8P5Jmghg9w03gInfuHadNAgN0y9gwYuzbrIGPE8iTB8G
aYBvQ0jM35xkneBLNF++oC9hrBfhQP+kWO+zXmLRDyga5Kwr3Ds0CLVk5eG9f235t45/vX/d9Sok
D1QJHEmuOM6UX8rSdNT7VJY92dj9aReKuM67/2lE1qgx+lvH74FooXuZnpGXZTn3uCtAn52xDonk
PUxa1Y/Dr8r//QfGsR6ZcAQSzgcH8kVDyytL9VmsQmTilyztfc6hIresGlgx86LbKTCM0PEIegHW
Xcb1IFypvTViv24wZCE58R8hcp76ET/FN8PxJvMTrkuUxMC5Vx4R+0SApefESYTtyMNt+cWf2C++
ZKetjfg/GlhZqW/LGehMvahOipvbLX+d6kjkQWxDsAGUmoYfOYosiW/4nk7/TEMQwOHHorH+R3BU
rvWUv4phRv64OVfNKTZqDn/y/yR1uURURs0nxGpt0UZh+f1Fb43uSuaeqzKq/8B9U09xR16KWowp
RU8xmxeadHVEa+DqmZYbvIGsORmVoxY1p+V3yMmHpIo4iGDeBdc52/sT85IIxcnMRCsSgADvrDdK
zgw/dHPRhGysNYeOBqo3+CSFAVs+tVrE0ugEQHoa71e/jUEzpWNSopl3M7Vkbeukh1k0XnpDiWtt
nP6y5GG+B07tB7KHDyJiNEsiB78XVdA+Lk1Pc3vZi27WOfqqEUVufeaWCpfD6U/2EAD8jqCQ7HYv
f3SLqAXr0yzXVuc3wYxC3NKT7epvObhC1WGte7lFJ5RPj45l3I9euAt7LEfELuMJhFVeqagQV9C0
+zm8J+AFLTvJosejiBZmLOqj0qx51iSCqLCf8x+Y++oYAhbP7veUzgA4pMA97M83YZf874DUaj7l
WanjZTchBU0eCkZT4sKsYwHlZXlTJrCGPM9WqkdDjUUe+GCoQJ9CUGVXXBUFwZezHYyxzApO8jIi
UpS8leWOmpnDTCqe1EoKdD4TL0/DkymQ6g5NzymvZafO2piR7YlUIPjknoYT8tHR8FHZLu2VDGOA
mH4ykF/eYQbzz05HFOYxCFEezSSxaxfuGHFe9ep1OXTxHKVui5QevL7bKoZzvIt0ezPEPLp5XnC4
/M85ULasB37+MaOwtTwBgm/8uKOBtEZ7AsPSm0I2hwfvlUk3Nlo58Z53UuA5G3/28l/+dB+Ij8CN
dvq10IRiK6x9TAbnQPQjGg7a9HfPdGUv/uo1fwNPZWA/ST9qQAIb2wARS4Bc0I/oQTjqWJKI2olV
+DXvJQ6WlhFd7rsfw9SZQCkc8xqdEL2DTcYCmguM8Yz7Gr87WMhK7/cTRmzksJDdVkOoRacpS9VF
We77w10YurMKetarwuo25bfvg872xSX8M+Ys9QmWeLiFYUqwCB1HRB6bY8f695eFnM37MuUxgPL5
YAZKIMAGy1lzOf5eY6d8lyqFV0HvzPXo0NXeaOVAVna1HFzWirruVVJEO84xdJGNGwlmL9xFSGUL
MC5cydT3nhwQgO6UtNacAGkPKgFy+M6y6PiGEDmfX7eK5FUXgz/g3p4SoyFexs2K9jzICD4itNIi
oZT5vchfuY0tWi9JbiE2vrDMtqxEIasH+Wx2a+Y4gezLz5zOCbk4XkA+AGgl53bzZczyMZzMa9l2
/YLoeoTGnNwYSOS8XjxqgOFf4nEUsOrQz2/eUmMO+CWptmjwQKz8NP+ECOb8gZH6iHNI0j8aDujm
32+RUNBvkk2sac+TAD13gTiI/HVXjRMNQYUr4iV1KvXIZUk23dj2YWNgKHaWtTWuWNcTrBCYHu+Z
axyZ5+1Gp8B4G546ZDy8EG4x0sfqZvpEM1Hbr6PHnmO8mKPfdCHWyKBuvF+mWLIMi0b69MWnSix+
KmlPwskXKqM4vVXMdLZDR/tiMTL/bYAM7aXyPVjFhUUueJz2vKRKs8M+VfWkE6rrfa/z8E20JSDj
B/2oxHcFyng+xJlbjY2Cp6NpIlr3JULk5PLAobhqlmGDWyrOI6TQ5lY9jiW+bm8Kn7liuj2RLrhM
bMiorBS6AKJuq6dEDjjb0bAIFXu7lMNjlIaZ7FaD6MrZb1bzaONYeJ2sYb9ESiWrds/Tr3OXXf8U
TScT0SKAKvqZx3JrE2mbZXdfdbViwzrE9Iv2Q1SMouEv5xuBZDc55rMsDW0o8jeRpm8ZT7TpTIv9
fF0VCUK24KKRtUYOxny2b5ZBwnpXXbSh0guJI8r2xJiUH8XhHfNZavMhwB0b8h2vlNU5KjDCfPMZ
xPkp0GZXA+z5eP1bnyZFkyfWtGlVJrKMnZTcbG5/HGsf5OzF1pZTMCHphDCGNutPJ+jIeHYJ+osl
NoGp0mk5gmJfkSURF5KekutphtAn+lNa3z7GxqOZ800moytAp33kWcb3dnl0Tuk8gvhvmEItAQqD
ptQ516euCvh2eFyGJJhnKCtvmFGhZlYFdKEcGxDCETu1R5s84RtpJVtwp6Mydu5vkpIdk3O+IMlW
sZq1y0R3rL3LyECx05zTFG6FI/VH459fRf9VaMpKxSZKZV8aUjRmQ4WQjrnqVQ3ye/29aJk0SKtQ
GMDGnEhZBsCOCsT9vFFtgdShs2E5yecSoBM4ZzAKcLcfCrEU6I3C4ODsqcR5zBostxUUzRW0qcdA
znnGxkxbWPc6qBy7o1NYyX0SxXs4/hAGGij4WEZ9WSLs/cP0MigQmPbESz8sxHxoCn554UaTQjo3
oAUz3eQHjLSpHCW6FszgQ1ysEK9OaLoZ4gfL4cG7eF7AP0ThJe/IuacLKPGsIsJzObtBXqiARifj
XVahIBMcKpspq1M1XN5oxndaAkvWm7O+/uy2XkEAvc5ckDAJne5t0FQlBVaFnbf518xlYJuw3jiJ
wcX1jJJzlfCpkMHiiPBL3zapGuN1wp262Ad5+DB64Ozo5RLNIEfs72SATqVKFKDLOP695tujayP2
i+lA+TDoEQnHJRfrNVoDqlRaQfwKI7y3Laz79o7hR3/XfkAYlqhjyCHzK3bCIIjApVXDI2juqSyd
3YOd0ZBSVyuJClHBkyQLt2sdQFOuXKc9bdu5dkUq5u/LZQn58n6WdLHbTJkevRe0xjRke8pFVgcS
Ekxjtxja5AfDESYQ/srdwclw2PvuPpyPbTy3y7wL+qJSslg/CElShe0pV86CtFNXNNzD+jYeL9PN
/8/atpbeDx+M5v/Hrog/cQWzpvke4iwBOESM2Erj/SmzpkGJsWR3m65CS9LpvBmN0Px+FRAybP7F
scZDpan60l8X2YIvtZdn6OU1+xrcRId01a4Ra1KPFLhmhqAiYMdlm5qpgb0KPFTFFP/6qAgz0+vK
DAHwkDUlOYqVzVEy5MZWJ1rc9sQJccEA0FOPN+OhM89EVKAhXn+S73/YqOsu/TgUhz0Ga881aSLS
e608/3wTCO3rOeuItS+IKKznDKEJmqc5FSToFHgt1pc3qf27v1UCOqxGhZsDGzSQYWIWidCpkkH8
D1wpyTfIuvLUhCFnHzxbQvansa+qO6BvVMFUV3AzP1msu9mPW7gQX86rlR8QFIIn2noDndDn69r7
Jyab+e1ecgffEOMzWX5v5V635N++UWUN35X4UtMKZ8Bo21RZr/negmdPByec4ClfVJwCAd8J7Jeq
RExydSkhKXc2mii1DscQ6ygROxMi4Fd6sBhtvCEo8JJ/I8K6f+7cnDogq+Vu1/srY2AdXwqXkXMA
a6RPbuaF/zkUKRJNJfHdBTE2W7ehiuVk1xnEp8DVU/3osdftYquoPTZqfzgYE5VvP8v+BYRswp1L
cT8Zvrqse0XKGh+SUTrRvGr6Fw3cUqXSg+GKIiHXpamFqQJHfH+PPRXmhTvSTgXh2/tcjtXVCsG2
XImP055alY+XigVIYOQwSCJ7tvX1J+nUMUI9fOxobuHHfgw3hp6jZJ6F0J8smjgXFnqnGpe7L02O
QQCdDLCXH/aFxXSyUoeizpbJc9cpOIg1YMvGj3OCihKpFnguM8oB0QVukU0chIeWf1tk2eMHsv4p
6BD/P9srnuc5J3or60l4kp/RGDzEJ/CWe0BOXjVAk6dLDgkp3cAIe3RpJKQ2nOop4bev4YG4dE1K
cXTqugO62gQuG693mlXoB6I8TQSjYy1bcWpImB1cCgY7diT17GrMur75VA2uOuGscDWbU4NMN1Kw
8xZPTieYlCAn2p6K01/OmYbTBW8dZpoMGBw7FIC4yZE27k4vA+fEzPmdy9CuQ/zdZPexRg1bdXks
DrFkbkTbN0rlTyHjSWrKysbb/qXxbqCgjc2EAE5neTKuZf0ysY0CyokAIOYMwZjtscoy9f0Pi237
QS9pXSGmvvTtfGCBBgcNru/etEgT4g1U2S+CCIiddk+mbUGd/w4jM2MkHe/LNUEJFP2DnFEDFfAr
yRt0lUZXUtBdaG3aQcUQJEw+n9gNDNXEsWZygDaTJYox9jaPxX9gg8mlo6IPJEkBULR8eqPY8jMk
jxrIBrPSY/7VYCxZbShG5GEZUanEUALlrS30CrJ6AKk9EvjVxez2BkoI5MMDNAynrTxqvSNem74v
wE6ws/j/KX9PwPOEoSJdVKzcuKkIvMiK2xFrqKcbVxvkLZeJnBrxHvsWWrrrQYRRDwbALfizGggD
94v40OF9PjCIzH33sindfM7UbAjRt0iqs+YcTdyiOfUxc3R2xAT+r4BU7OqVxSN4Nn5WAzKsOi1J
S3punEXG7AJyfLusAt/q9/47rRHGb7KhdQeMoP+aGudEuI5/5fIU9nVRtumCtbtB8b54SrhU4pi/
H+PLHwH41rmqZMxFjSP1usMiDaXMSqUTCi8y/CkKdM37Effh4EedU1L/XUTi2IUyZEbK/6dOpCg8
C6dPXRI2bekLYg7jFhHWEXORjzVioa+59aTP1H0Zck4Q6o4ZP+ktksb7We8zWIJnP+ennlaCkQJ5
EV9ioBRYUmvp6CDKxmG3ENoyjnaw+RiohCwRgVq4RacKkYL1RVlIv/4YYmgOctzWaWwUd7hpc+0h
pNE+zdFDlRhi1PsJvAflwd+ReFSLLj+58U7QJ9xlgHJVY8JYaZEwlQA5U2ucoXLqpP9WORPCOb3y
QlZfMWZgA1OOkJRF596wXaGjl8Uvyys6U4miVJbi1/PUavoiOo3IUgRxOG+01viiTnm2n/pQbLRU
gdItE6CCkw0ZW5JcdrzbeNPz8Hcno85CxL1D68kUWT6rslm/dIT83DznhxAQZDWTbzIV+zpQCzVQ
y6V3wjqJMJX1txU7OMXUWvL67Dc1SOFXookJXTVPMyJg3lZGUF28UvwZUI7KVD6DHUds3HQh0a0G
5KWNn2wbVzP/tSnF9cEvaDIAAdmjv+LpPldb7i4qnM+5olzL4r/7xZFT4H102h9Th57z/GZFGHtR
EMZlzgJbio78Ug5+n0iDz9NZsVHVC/JYvqtVm0Q0Ptr6NfQyqdMelMNU+1tqv816m8518baH1W18
cN4ZMiSq19jppj9wOxhAsHMWHly4SPypa9kVwd0lAqHrswPBFxN9ylT7gmt1NbOhEJLyolWQ2Giz
aavp6w8UQ4hLz65QmnEso9KT9iwZBepDui1nre92WdmeL23uWBCsuxDSypnkGKV+3eGzVl5pt8bH
4APVoPUUAlOUPxBkVwwBAqwSg8t4TVE8Yc/H3n9DWp7MREGDmWHZE2APDWYpwOVNDi4a55gk8XFN
F/TX+dbfXgbOP2zNADaAp4GVKyEZnagE2BQ3ydEZsNMQxOrDpgzoutkZ8unfjAYEhvmQdZXG7K3X
xd8fiapbMIqXL5n8k+OwfgkGioKDJz6fbPBk7r83k/cnkVCNwW5L2o0jIfJ7v8Vh8whgZFlJP5Gj
OH9UbJECyVLGn61DjLKNduinSpaa/ZGwjzu/8Mk2EhdFAz0zAwAlZ3Q5LOrHYCi9QxtIwIEQansC
5FkHw9D3Ttr2I5DF8/CvE+SwJNZ9TpXeLHPOOk+2wm8aGGsffhCAIIn8wW6PEfWjMzWfCw5vLhf7
auD4bGNr/eIVSMv5OsPMvmtYQtLVKcAVifCRYSZuJxJX/acDuB1arNjCjimnzPLT3gIfVsFcl7u5
BPWAOH/+YBhVZyotmQAhSzh9apWnFywcMxxEJn8iZIw7cmFCWVfIYaNpreIQ2msNNwWsL0K2zcf1
OwBhXymkH8ZQt8vRetjTRXWVCYGOKBJBy7kAUnQqlow3P4rDC/u38mTpS4VypCMsbFF1WhZ6h7fK
mB5iucViClER2WoM7U74Bhr9qIL8cpaZftyir6/aMKPwC67Ia3W6BpYgHkkydvkQvfWL01Nbet2z
BQFyG8ZEjZKhFDNfYOxfsp9TQOEZWOMiE1qjnJI4iz9GELLuvafuc5wI1K23wWTwuBYxtxbSbhha
yG+d1RxT8D00TIpEJ+ZBFBsXJF0pV67MbjmLwHZ0SQ1a/RkT/lrmKrX/r0/N+dF/3LPlyNa7Z07k
UTyZ8+8oBCakvwNovKRpwOS50espgCpDRo0nSLIH1EtUzS7HFXL5g7FIcTjFOWqJwtPGxhGUqWMF
U2NytVWihyeJw5BSuRpNRPp6DnMVLO3CmLtq6qyNeIz1hPCOk34jS9w4pF48ACUbuEMzCf12OEHK
E1drQ72CBD8bJYKX/cgokwTDTzKWwICNI6LTrmJsPbYrtovG1XF7sbcOCSkruReDEuJTRc7Aorwn
k1X68B2tci0jstaDei2I4f+AaKbKnAnFSYbTQUxCv9VnxyA+jgBqN1cUDiYweFTYWkxcCAk5K51f
+jkPjQdCBarHCBsAQMLVyEZpwGpKJspcCQr4hPtRkp5vnTGoVjuc3c4emzzvrNJ44SqYkZm7j7Ku
Sw7rwX74Qv8bauxBYaUJJWA2uDvGuFZhfVsILVORUsG7kHRQ0HvSaU53gHWDpQjA7/32JQs8tY2V
BGv2Na2r4xe1SHJE5hG0+5ckIfJO3Ykt6pEy7tiamGUoPPTmXf98dmAPS0uqBEuBbg6hQwNoS2oO
Ekg6Ns3mJ0vhT1JkioQ3xcC95tso0woVwrkFARWGBqF8dDL1OTsGYNcuNF0HlJ87EYWLYLrT4xWI
iFGLmP49vOWPZu2ahvuzvYouc1XHqhL/BzrwuJlBeMKnXrUG/6chriuKjV/5xVoUmiBqfIDbTY8k
uU41aBRZhkT9+yvHiC2DVQ0f8vsYLj1HQGx3RnOikZvt77Z6dcDT5jHGzPIFnKHnIE1fpSzWoqbF
Iw7WaRQinGdw/tH1CtqjLzhnn77ayxpvOc/uN0EaXGcs8W/ZEFlwwWVe/6+NTJDI6n473mAFugRQ
Onb90kG1WaxFDXfOzZGfyWSGY/zRMMklsY2yFl06lxtmGH9lQBO21dHbK6+Sk81OR15G3iad6nPa
SS1Qd4KMk39qkAJl1IQIcfJtRoPPWMyKGfe+iJXFFyr+j1+drpynK2BitMGdNctCjdzpIiedykwv
KoRqsBj0w7UFzBJdLK9jls4bKpAsUzNzXJ8e5I+UBZ1D82N39D+3RsG6AUG7cJe7Ip+gTIXrFf18
I+AKrjO8GSL/Nipo/HveYKpa7OiLnA76OdJ4NEIDHzPmSISq0bGd5bc2UND0mSRElpJZP4g9FmfS
Ll7tCtMm8gUUkKLcGLAC9C56l3n3TSNxm489dzSZloM/8y8rjHg6DB24QhCYqGB27ALJrjKjt9hZ
D37Xu3UAXgOURb9Y+/zRWq/LAxCxtQib2VqVkyPwQfBMux26H6oQN8HKPTy7DdqHoRGd47WvdGR1
yB9Oiv5rzWNnyjDVdm82Dwov2Otx01ijPh3v51hIIE7PjR9RyZ0DLO7I8xxIHowKrr2/6NNdtKG3
7p/Vyne4TRE9RaPYmVhwuWj86xJrQaXKByZGEQ3OfyiuiS+T027p5znN2PAoTBpET4/xeDnFiyQQ
WmJ+eDCfIvrP5ozJ9E6h8q8mz929WYmq1AhQOjguSFATfZo1y3yCoFExRtl8vCRRxfE2WoRYxoxO
Kz6wAzRkl7i8hUlgzZFTs3u1MiPg+9rCtgMMzZBdZvBa6ONSV2ouqJfy9khkd/F+jR7KhvYvMlAh
H5OwVcNrAkgrOB2jeh+XGw86G/AsUo9Bnyjv8O/Knndt5gDnrpLPVcMWZzn90kFUREoVvJCiKUw+
3BXHV6J8wq6TV6/hx+7pLVTQvGPYfWkA1/mwgLVgBdVJkUKecCKo/9MitykpkQMiRX4FvqhuvvoT
t1bFnP8DhDuahL5EiC7Q7NRnEug/G5lEu5kM9a5vNAjzVOvzZVcp81oMmwwMnJJD8AsFT+GxNiwa
eHLHy0LP2I9tMbBmSJB2Iw8e5JVyzbLZ+lCAaBMBq/fhAlDYMXCGmesepNLJj6SLLALwgEplL/WN
bN9G3bbVteszgMuvrF2rL/eJrOAwbQsk7Tn0NXgyrp6y09875UlWKaqSxGECVYs4iavXK0vCS3a3
MrLUKfcC04YLN+1G2BU5GXARNr0XkXL3RQXdgk0DEgk6mt1+gQ6NJTbRDREATkNns2HIMbg6JiUF
mQoQv3kG+uroHf31V0wHeLeY2VQ9cEhXvNjZ2/IiX0M8MGkVrg2qwxMkuzXP4SGCGZEQfLkohq2X
xJGg+9LNuBrg5YUXq7tyv4CziQiUWrKXFukacO0xfqO7M9wHfCV4dShP0w1tZLNJE6NJQT3VC62w
s/eSKvawSzVAw5w/ldy+pcRdSlSbhnCM5gPLh7QbKuUXrwDJ1b1eN3g/YhFmB0o9LV8wmdGDYDDz
O/e3e+5YmOkbDOc2sr3H2DL2MYFB3El9X+lUEGWi9aWjpf9CXjYXwny8gkWpBBkB2jST+c1ueDsW
VKMHNljkK0p1AVYWJOja7t86akAv3+g9m/ouXz0nA5wt0B8MDhpuKiJ/Bw8MhvSqCp3kj64tYooG
IwR7fDhjb4jGztSnUY8PlQ3qcbtmvQFpHLiTZQ6i223GyDgDe1FEQAozxRsXHw6FzWvr2hgoqzIz
16MQZiQWJ5B/FF26yUbKliuVZooaQioLF7NSfr5lgPl7/XF/yczeVbsVNucXx7QKuoAvuKmlhh0W
j/I5dgrB3agZA91MkpmGIIkmpHeYOhirg0AmSDGqhXtKJ14jKfR2gcnNh63CG7VBBzKe0hm9QfOh
KhuN0Ju3XXLwPIk/yvijIFBw8CcubpzL0q5fcFRsNr7F2E37oXDD/TE8Va9piGnJBmq5ypd7ZJT5
XaIQ59qOyG6Kvi4LCMSBGtVHtxFpxxU2RRJbUU8296Al6EAUGGCPvo9zp/siJl5VMDYIJSh7/Y0D
nVEF/Aj4McsVXJFZTDRR0f/oMI8nLP1WcXqIDPtYB0Hkdq6TCvsPTL4u+53DYHwjn/TQuROTfD0l
Zmz1MULvnz6IuPB6zHmfnYW0YeVKDi06BMUcl87U0IzzBa3SL7Y1Fx7eurmwo/twvUKUqI2CIi5X
CuJfrIJ8kKzSytlbYqiCsKJxtZvVJopOh14saqwuzQMjeRt7S4amEHUnywOKw+GtyeGNgbqL3wFv
7ZNYExMiTHEAPrxZLKpCOoPUPNLMC8MC15/DgtU5VjKsOIfVM5fikFAXJRId0oXn3Q0TFAX0dVtr
mbiaWPQNFJUSdzEnMf8ZStNTkduSaMeRBqw9riSwxr9TYK66z1EJNYFWlUIiKjChJlVFE/aD3x+N
/HfgZkwTDvuKmHe5lbyrv9gu8n2jEUEfXasxp7Yb7fTZUF+t8ydkjREevqrLh7fNIxbynXCfzIx0
z7yeZeb8eh1CA4wkPZ8s++CiqUeTfoOQ/kMCCIYdyDTEqqKyDTd+cf3CmVCjspGpN48eSDBHZH7a
jnwEDjaGqLbi1DeuEbnmMEVjEh1ZBj/HDP/BS/a9y1ol6dEBaq+mcI/mDJZMOjX0Bhz2WLwy9v3P
HzvEj8rsKWgvF/eTvVr+q2R27qfkfMLCx+VbDvRWLgB7r7++rVRmTxyvfsdWj0kAEUkQeuw8HlP9
aqYe6Obz8tFUkvoK5LGvksd2zOt+pgD3XIR4hgNa291pdSEbYjVVKRZ99wl0hTQOxOqKmNoNhT/N
OO5KGIBzdwb1sU9WraN3M9qNNcgs0K1xdEQu8OIBOQSIfnm/fnjdxrDun82nZn1jI02HlNE/29S9
v5b4hGY6Yhp/XRAkqkPZTpPYRstBi1lgVlcdu62Wa0sV38Jo2mGL4WWNSZVc22l05euyhpCkc/qt
gHjm5BI6Tjmg+eQu0JlES73aDKRRMoWYRdEWtInQGMtQngLDo3w89DyZkbnyESWz67c3IFhmo7WW
j3QWEhdimkB6ncgq2dwt7/eQyplvYnp2Ae3brxFy/wJGESmJlDboIsRj8xINI2wq+/8u3Hj86CSm
oJbajmWS2MrBgGCWtiuNtetATBDneHL9b1gQHcHGVm9iTsIrOeiH4tvOYhOSiYt6XgJf9ZNI7SBk
G0vy14BXQhxr5LsW0E/tFLzZO4fes3VDR8a21s0ejX3MOg16XkIUWqXSMb0nOTxK4IwMbB8s03vD
y51bjuQ+apQQMsL5AHksYjkDnXrubn4/vDFMSuaZXXquy6S/sPkFei2kgdab1A/qyzlWHFm2rLoK
ASewkFuNFsrwLYAejB/pi+d978DmFsmiCmlRKR1bw1SQltGBr00hA+KPknQvpNgJZPHQFXM5raS/
dAf44at7qhYIxqGNYYtadF6D0XmWZ+mRqkLvf5QYOybuUR5/N0jvoLs2KXgX+U6UjQgnijkcnj1A
/Qut+HvbvqtPxx7EjoepaDlqotilW7GEROA9nHnljSLkJTKIMUbwbfYmlvFi5TCySJXBjheyA3/Y
hz6ZaoOpM90yFApEb1yNMBU4XJkSTBiEtnQE+0B0mSeTFVAigEhDbfgHsrjpARhRFmXpuG31EpP8
Churkb/qJow933Hexp0zO/0HfxOMnYFuEx4HvJeP1XxjwfyjTZlXBZF5eeALXOrMoLNqTjUNZhn7
w7l2KZPW9gqJHoGOBJELH14cO1+bjwElx5sR97wPmIs9v0lHlq0v96Ukw2rxduEOBcVV3yeiOnio
pdtN43uoxWahtPdp/K7Zuu4Rosm9GFyYdpRieMJqlGZCNy4DnvKsX+9sl2ZlcIj1whEp4tWwAKFx
2FtkYuZq2PeYjI28LzlBY39hBO5AhrdQShyIhuqqbPcgF5oxP2oUa5DIhAbDjHblb6VCqf5P8LG3
aw2oSPwki701uIt82mvRdgckvkU7YM27pxvWvLwvmTSr19VMLBWBFVpXj+U1439JteT6r22zMZvY
LTSh0aaytyZS6LEBWgP8prQN3fe2pfqx4TxPYM8cTTF5qovRcoaWVQnNUNrHFKNDXrOPeu+mirB4
HTKEJb+uQ/Zs873XNARRILmTYg8FViPXIm9YJnfrHqV92OqAM9kM3lPWBJcSoejn8n8rylO+oP19
Hg4tuG1qVTa9Gf6wP5yFLiV0YFBQu5AhogKzLkHdph0Pd3UvOZw/hpZPv6DsEl5mafSQP5r3C4Oo
gYsb2Vtfbng/pUgpLihXtZGoDCe1xt38u/+3wb6qxrLZ1qURzhn9/d5qkpxWwzj12Fd4mdDtbpmw
KIy3+GgH6TBsZT9OtmS+owVFVdpKDs9VYPzb3V9QaEVhEYc+3QJOZgGTTrtJ5AS70S1cQBpGfL3m
9lLBiwAPUCFu1dkTb0eTH+hMvE9JHDRpaNCSqu+fGUeYV6dIt5PY/cdZ0gGqSBIZDsgbhGX8m2+T
9I/9RDo80lAHxIKds2SXpdvCbBMQcoCggzgZ/ZCnrb0ZBf5BM15PK+I4Bhzp33iIHxCNEVkXX10s
p4CqIcOWSBf/l076R1OLuIONaeGz7R8+nu0X0UOvtWmxnyhFtLjjl4yiX045eAwBJtupjLDICowE
1ZFqyKN3pfU24j6AxmoxXPJy1iUdVSvPz4t5+KWoGePkagIkIbCGcrXcrJiPAifUX6y9ACNsigBV
9W199uXiapLRzYw/oQuxKt4lp5Zy8CacLcxMGPH6q9QptrcdnYmfrof9m9DHJLetvjMCPlMwQvMi
QuVSVbpMg6pZOLmJRa5FnJIH6f7oWCMoANcmJ65lPMANIo2V3pQb+hbUg/HqAxxgjIy0QbkSB0zc
9lltCkcjS1mVSgNq2ceowS2RBiIsI2z5Jz9Rl8uo1FlcrP+7r86f8JwS58sngZk6yHRLwfVOI2wx
tzhbgPGf1kq4fP8lVN3xESnl1ztBUBmzBn2eXI0PWyE6Lz5go5bHzdubYsKIGCD5TzQf7Jjq+yUF
h3ecrDfXzPnmffREiSvLGfSvPr0flowThVxBsd1v5G4hRMKWcu5G12T3lWRw3h/aoTjvRyHd+LsO
PeuCskGVBRd8vRIgIkzuIk9AyoY1lJhipaJ2pCh54odk1OJfhWfdMnA6qARZGAQk92oc9/WcKv+t
EWKzKlPYN8ORxe4QzwKFlkGQgdJ9XdiRJlpLkUE7lH43loJuNNZMoxg297w6ZbGm9Vz4rPDV6Bon
+YbOE0JKuJA/xXDn9zc0cdHk8k40q18tZiTigRTZdfjJ/KYwdtEU6ufAwmw0ZKYUmXFJA7TGj4tM
V2gsEO6AkwVRXRi5cSsARQqa86pxZ3oybjCWxK3u3v9qVTIJH4yZ4AKAHydjb9XwYDu0+dENabm/
Uo8zy646uJqgUBizrHI0RUe6ZcEpiroc7sH8XWD5+lSaXOseAgpJzkuruK1v6UajwPa/lRd1MR5r
WLob3k40TD8Fil8/jrzl+qG7KuU9bUcm27e3iMgdz7UXcsYj48UOtuXYshUbCNQ9pOTJl5UqBC1a
3X7OfmSBKSbvgRIOOdtbBgWVHTjzcZGYvsIKfU1vNot6HRczI5ITy0JQDNI7JismyJ7w1HYxq+Vg
dNWAgWmD4be7vUnXPTdsUx9M3Hl+uMDeQIdeajMnrZGV1JMZ12FPaFvYgaESZDBBgEZKHKFRJ4uC
C7iUo4NZ873bxqnIHk6PCJguPtnt/naaau+xXL2/PT21KR9nRxovM2/Aima2RUmNd/IlOOMVEsCw
q2MdR8NLZ2JQRB847DNP9kO+7X2NKOiCnOc7t1adzdXKt3DlNdWykebr9ceRVd8GXNgUGlnA2OF3
5tEo23c73laqq14zgGeEZfcrp6cJ4tffDIWT7rLIhjaAxLiq49ue/bwojXfx+zGWqze5Jr8jTsSn
PK/eLRsFDm3wgJualQifgT5njFPc9WADdh1I9/7FMpwxk/J2MzicubPnF3slTQPhZE/qaByzdTWp
ceUZKLabaO2rrepXWuadiXgMMw0kC9n8HAzeaRyIkKMFxsoeMQUJgjGtJG41Veb5LJYGdoA7hFD1
dUsO97jEmkVF1V6R8iLcNsIo+ReOnnS9u/iXB+Or3sMIPCkV5E1+jYGaBUA524nlLMxLrv1JDAB2
pBIo6ldGzGGrGGTqW3V9KlH5f8n3ISR7OmkJHJBXOi8Sw9Hoxk7QhVBkEc2MxqxVg4ifX2b4Ohf5
DOiS0c+i4w92yOMhefUwxKXaHefhexMNO5iKv/kCnJ1r6nj9x/oIl8gj14lqk8OQaP5mXn495m+8
E225Asi2Cx1/8CCztQ1Yth4R3+N3sTV94NtHHDuzrdTVvIXOdyeEjqm1VoFf2g2xI17ttHS5m+RI
Pxl3xM/Pd7W28Otm6FMr5J8L6MdtqgOsmt3Ltfs73oKmT+WDrVeRZv6xrs2+Avp51gG25j5rionI
Biq1UbVthA8biYMfviyOWxr9OtEOCSyPjw3isLZy173nK9LsyiPtvVEp8jljavBnfbogLE4ki7OT
OmpB64HLkNMk0Mp2lVQdARxu2sMVITXBoReb8nuY0Hei5EQhlEB1SzM721bPHXp14bhSlx7sdsL4
cA2fqI9nDi0iw4GrI+IE9XWij9U0gheBVXmEtpZhutspNDXJgw3C8UOPiuxL0ftOCAMhx+EvislP
9wxWBYv1JGT6K42xgXNl7/drvoUvh6pxQDXhF5Y8bhPJARmrOS9Cgg4wg0dE8mMcYZRhZZDgAsQ7
72jQo43TOfhOjCbh0as7mdc+v7jtU3Odv3IhD1ZqakIGLryhNoIKyJeh6kgVy39ARtrrj9BStkzo
OIuRPhubxMy4iYw59XRR2DHv5B/8wF3vS263Jw4Kkq8hB8VVbPOdBTa7X3XQaorWaXMO0bDunK2Q
h//FojbojUZjv3ekW1fmIcHatqtnye+nWZ5zfmpJNQDGxB+8hgBo82M0Ng09bJhtOv8fFk4HDdQ0
9+ENvS6Xdu19AyZxKozpnOstO6LvBiM/drZNVheMnGX8Th5QwdvAlMTTAsEVmQAmKc3DKFsk/P3/
srbF6Akc357BUQeNq8/+vM6XTvm3CfJHI5bQEZXq3QAHIfpgVhfh/5cL0t+9bANJWTD3IoqESL33
yZwbQj+ofM8LIubA9kPLGNqAhlJg64sexK5WGk9V5TNI0b8/4YulRrmz4LcPw2EjHESZdXbSgJEb
dVt4V/KGWEOsmDQMRZC3U3aCmcGO9MeC3ZfM/QvD+9xzOsnGeLH5xM2AmYH/wSOi420y42x8axy+
OOpkzvUU+LY2Iz5MiU7OVUw/RdtSL0iT3mmVv0K9BcgcemK+BYqcjiOkAACjtmyhB1qAeWsIUhyV
2Y7BbK4VyL9MyVifLKh6dtQ396aPxpMjgpLA2h2U0vE2G6dm6GjGzemiTl8N2DGpLlM4MtVwQycJ
6CLKAStqf97lgW1KtzegxRPfDDnGhqVC0XSOkkdBu06LfPqUWCwrFN8Go2FL4rdQXhhtPAgP8dxS
7ptgauzzWRXL+p76RXyyQIAVND+7EpdUNu+Ggv+KTE2tGcRnaLiWlyobSX4YAlRjWJWobWQsSxIs
htywxS0jECLqQxggAeiRKVmWBOfn7R8vEqKdaHBy4ELsal6EV89Gl1CUjgYODyY0B0aDEO/X7J88
3NNZiUf4D1x7U4Q7jzi27ri69682ck8VyyoN7i0ucVTbvdQBxv4lPUAk2hXevHUiW0+Ed2QAgT6U
vEidov8xRf4bq6BYZcStklaLJNkLmMf704Pgpo4RVYTOK6bjNHM04NeQBS4v7ynbVUKf0KF72y0D
1VchsqEsI0aZcT/gfGF+9igiQkVsVQ640M2DTjQ2Xihiqev3PfpDCzz/jxLg2G46s8iXcEbmKh2B
3TBeHXEkKRpWMm4S/CvtZNIl7wliSdrFKQzCaLIETn0kVPhyUzMMgPCOKn3LkSD6yfxGU0C+v4Yb
yTRyAZ7Gb+1bq8HJVcXNNLIhtkapKRI46qMF0hkXFkrUfLLdRfAM1IfLT5AL6aFCG/40uqEMeJXJ
7C8eIRkzap7ZEvIuBjyx0GSGbRsVrfPJkxo+GXBlR1zS94XRvPLjgW5kXNSVo6KWAC49p6VbEWhE
KPsF8cfowRDAlMBBNJpXpS/WRPhVjfGCjEkCN68HfoLb/m1oKvulC2cq/PTiGqGv8LF0yW0bznnF
kUPF71lLePAwoTQk9xRQcz5ZdjVTCniF90Uyp61/lz4zECZsSVxhF8RnvpXPY4dPt2gl+kTI3dnn
vxjEehy2Y+MaeQLQWNA5EATVIL0LwcMmwQgqEBYVhidkg76TKrBjjgdJK69wWc+5xOETckiV5c25
smwIwZqBHNAWLPf8qX5hI6SO/B5gcqMZojzaKVLoC3ZBTkPvDv8ezFYzK7J/14YpGJah+xegrWhf
Tp9pY90vt+pcaTx//90HvAD/MKfpDOvJA/9FvLAQabvQODrV0K8cD2ril0/ijN9t2moUtaXyYVg8
hMyXreGG4/2EPIEcSy4CGXwFLHbIkaEqaO265SQKPjNf4P/C5o+fOezs8nfgSNRe/pEryN5AWDAr
0DvKuzO6IWdAr9X8CWQttcgGnGFEPNIPHrq9JN89ohDIb7N85mMjGEOmuejd4re4IrKeb5KyVOdg
3y7UJB+9nDaKz8vl/zPQjMvAXIYVZP/2UZrvdmMr/1UJ1Z5r3RGUMMBOfESlIdKFlrMdBkqqMJ8X
LFONURA5l9qCjzjLOKI9a50uebDJ0q3DytlTp4NtTWbqSnJCgAEuJvqyVcvfSCOi4IgNFg9JOb/G
PFNMSw2oxrRhTEpulK+EAG8NWspJMZXBCJX8qxdd2nrbNwJZwRT6pFlJ8IIZIxDoj7rN+TItEa+Y
uaH6AU9tOcLe9hHsRXWm9h4yyDHKuQFJv6Pur7NLDkzlfcTIKWCBXVd+BsfVIZ381PZKoX1e9WLk
sOtKVdIIUJYcDAgWEOWwlOvB0r+7+oVTvS8+pjWqJ33D/SvAo+B+SjZjBFrcQ0VP3LWw/eChPz0x
Ef21JCXENd+1tkJabSbn+mZ5kbxnLwVUOXArCLpqPO2DOhpBPc0T5/3fcdkdN6Jd1kN3f8hWGVhY
OZFM893sE8YDkwyAchIwd55MSUMxbW4ZKfEkEeUeRwRK4ITSOPjNtJPcf4oZ7j138nYYVRuowMxk
HNbeBMAnNzL4w1byMSSgZ0jlxw/h0N7lSP1DnxcOklKI3vUrCah35xeDqB9CrlSezcKuRAc2xmWO
IbfSADQ+q/xhByAvO/0rtwOpMMChM4aYL/ZK/bcb9Qbei0tp11zcL9d1DOre0GiSigEqGoh6X5fA
cVYKW0jYXLRJXBcibraYwapl8G85iVjO5k6h10bGSLi/PmjE4IhCC3nAOeby7JeGuB5yQH+IV6Oe
7FSdMiZ8IdLV/gitqp3QK05EV26M/ve1yOQ2dcwlD/i29IDIWMIkVuxu+K1OdwN9ZwTPz9FVaAFL
2wp/HUzuhuNR/mov426R6aEJ6bVeM7FaXe9u+w9P8rkuEckz7IUFVUWUjCVCn3RybHlHeSWq7vOX
4LuK59Qri0h6kL4UvuWHpA0bH0Vw5Yoaibz8mZalUW+ClRG9hZJmSX5aMJnvspsp7XBZgUksfKnB
2vZu1VnqF/q0Fnhzmg4WVEPAeGDk1TbFH+AeE0M0DYYL1VTUjxotsmFN7+vla6IsIbF2CQWo+45E
6y6PqJy9Nre9zGBZiNOHAv8cQ/2ip5DKhFtnodkZBe5JFBwAEoa7RbMygRfjVHG876avI/8yedF/
yPsVFUQUiIqCNGVhAXjQEq9bSWuA50G/x/BxOsQWfZED00/0mfDlQVXb/jQCNJasCZ/NPyGGXfIu
cTAzwTPo5Hp8gUfTZna0i8Mz1pLNoxLxpvGxT96Qad28ZUzhiliIW22wx0xo5WRgRvV/K3hX0sq6
0K6a9u6RAgMjUiHwOE10c8l99nYmJ0VXbDOpdFDDm17kAJ0jDeF8Q1xniownlqkBAFtGsvpqOmXj
3qMn9bYZ6QUIoDqS+353p08WLC1+6S5oc61XnQH41gTZmX7nRleHRV49EJQXfW07MFb6dGCp6/pg
NPBkHCqNtGzo9lZ/MVbBV008bpS5+00C7LI+BJEzXYkJkOetoMPL9JrOYsEdUYIWxZ/fjrRJ9EXS
2mM+dGjdinjdKvSoueuZjczrXEG+PCC+os96F6ybokPmDvOY/m4r4vFR0IXx3rj9HTq+JfKIYxm+
gf3lG6eEsosa5ZTzdAyf/hPJVfhHcqszdI/oraiCczbmyhEbbioifxyaB6P3ErxdlK+QcGPP+Pi+
91zv6G0V+IsZ/ziOznzUGTlWQnFWQy4IBRi7QmMitTQd2qcxig43wjd71FYqwdlYffYZPGw6jWu5
2a9F0ZAEMT6ZGJyLgdTyN8XPE8JxJEmKRCNYZzXqoYsM7YBeR7HWA++hMWqKz8LX+ZDaHIWVwpkI
RGQlmMditsd+KObL0YNpMWP/Ow4A3SN5jydOY5ndI085xW0B+6GgFYY2Ufws4rOEfo6eQDYmWfbo
PbDT6MhfZbpSUlwskyL1PrkzR4wEyY9Tng8uSsi4ycBzKoBllAWIUldvTdDParcO/x+AnEEB1n5+
9mpFoj/feWr51wXkEcbbDNdciGA2md98O0M1/sNV3TOSbE/Yq2RYayRQMJRlnAWNG5alODnO88pv
oGbIxvBE5GcxnabYhR1CWRXasYwGpnXW1cwK6+075fkBy55cPHQwzu2uL5KridZlwft2PjIj4PSk
fHGn4HW0JK0gWm+CSJ3W9M4FhUGGYBw5/DNq7OIKhdMH5b3n8IatCSrmNmrBk+gE8SZnCLJ/XYsx
y3SrDsqA/uHJCEgPbztm7qszsqo7Dxw3W1h3m26yiWQuiF+pXWBolI/CEkd4njJdZGsgRs6YrRrn
EbQgkJmJMALRLcQpKk4o6SOh0wg9kZOS6s+QsQdxAcf6Q1S1Z3oykKV2QCIh7ynZSHWoFQ6p1ycJ
4nM6OstKzvxA9IUlBVd1vg3qZbu/U6OoD/htqPahyx9AG2kcEC3uR58nIJHiX9qZaahlimapKf7l
SGLBC4zVFcP+W8XoTYRqdGQWeiOkUpffWrA9cADneXQFId7zvyVKWDgXkGT6joBBRn1ZWqraxnhu
KL9jHbIp/FvRf9eRNR/57rL/TbUegGW2y+FTC+JEYjImAVb5EKCyI4LDRrp6HsNiGVxndVpRv7nL
A8bR1I2dqeR2aif5t41SZBj+gTGUwcLrqnLg4FNOVYMRAOk7otamhWxYkD0nrKVM4jxB8XoZKvk7
Wag8m4d51GsMD0o1qDMS7XEULrF33U/qH1Asl1Z7VvzsnBJzU/HVj7akqZkDbRw1oO+wxLK+v6Ui
LhytFRggotoMcTJHJ3HppfqWbyl+gx85bcXBSrHnkBQdI7VCKoxwJdz6vTWytffyIB8XBzkYNwvy
0IhWAUO/wAZ2Mh4I60qY7vpwyiKwDpo+91SxpqcfS5Ht4zEdCfoTH9UERSz4LvsiX+c2jbXDnTJV
mQR12/bY+56yeUmlyh2ciu8i1Iw5/0kLUUghzBZdwn5EWFsLbJtJ23McEzxGRS6pbofXvupviHEc
EoyGAqBm6+peE2Pobq7iDfP+iB+d3MZ+gzeEu31j6Hk/UJ3CoiXRnlDcMFaka+xEszSBtvPoAKnD
/2k74y0rg6+29v0HeF/BqrnrbSwUyz85troMSTAseBm0RYmKoiAPn54DXlGDWc1Bce0Mk+9yBNYk
V+hWq4jkHuf/4nnF+tSv2zFzvBoRRp8E7iDD620VxvMUWJOn+P3dEzwytAG1p6Swbc669bjzhzLv
FHDzCtYkPrdczzWJzJqsLaFkIEG+fWlBI/QTQAcPJ89t37xIVYA7Dj5dJpjayU2Ti6TdPTph9ddT
WNKjCHZtS277cHNLjt6a6hYsbqmWXGkbhCNinxvRmBE9bx5utI6W5OQhnTPdwpUVaURju7ecS1m3
nJ2A2KJNbj0UJB5eYPJgidIQeTmhVmB06LUte8iRK3Umtk9mYkfFD75JLg6BL4hk+BldMsdd2hYB
aHmGKZgUsyXYLJx/hMHUV3bytwouR8ZAL6Hy2jSKNtPlwgu9Io7+IHPMQTTI6EA0V19UGT/i6rNq
bLZCYhFCS20gbvuZwihRO3TWwshTDGJZ9XO9TBU50NqAEJr3yqDVXIIC+xjPiECc4/MXL3NyzhUw
7/hJnJghmFrUVWyvxbbGKz4bT/HsgIoc+iqqtwtdqY1bgAXrLmWS1688YMJgbHNkbhlRuKcKXpRq
0iTNO0nM/yA0zewFwoyunvbhVIq3gGc/3Znr5asAa9AZOG0aqFg2sizAU9wo5fQACxPqtedWq6WO
N7lJXp07tIeFkAFgqeNAcRpmHcR5Zmc5nA9gzkBW4DlKwMHmF5lx+Lkk4SgyBUDFGQGGAl42xXoR
LXao7b5MqWMf4LBysFMKlUEEImCa5LIkIJkPw5vcb1C2lZz0aYHgU8KICJa42nMYOGlIIcYTZmjj
XX8dRex6Pft9oigzjLp+4Dks5jMGt8508NQIViKZB6ZhaGr86T/0iFFIxzyQBFoyOAKaVayhFXKa
XdICOs+cj7N9pnMkvQMuD92GXeZz4pYuLrdqJd3xrA3o511sHGVfx6KdT5EMH+zeAZOEFn421t/G
+uXqxhv98KerPa+RBdr5HeLPTXyFtP5BPWrnwnocq2WvCt3XS5irhm3u3TVKQK9/l1Afy/+dD3rm
I/pz+2SM8aFwXbQo4jCdcxwAhHnpn9F3BO50+As1NnTVaUp9dGw7mIYdFGOAN1KWhzlFW3lRgamC
XFhZah7tV8YN4zqNW1vqLfcUYeKjv++Pax1Q5UjWZAtrt4abqCZuc3FjwZ27ObN9yrWqRjqs5uYk
NKSRjAAO4m8ZxnfQgHWHCg95AzLAvMO/YK7A1Xmx09+w6yNi4Z8c21Gdbh/KQi+VF1ZNDFKtWhVE
IcNw/Mgy4HTm8XF5RCUZHvEHcgqJmJI5ynRcz/S2g0clCvsleLc+K1qvSIi58i7RWgRh+LlkMqXq
EFtwhjaUZBd9EZ24hZ3J++FeJhetyBpoGUUd1hjE/2ParRehpXWe0bVBSdYqFLI9YkOgLRsOSAYv
Uge6ZVxgjpf9cJDGGDrBpYTD8k5XwTGDbwpkaSDOqjfoB6I6AhPCmOnF1TjIHUroYq989iV308SR
VpjmU+5d5gSRUy4yoKE9zLYArIl81RJqDWCyuqdUTo1zZB179vNxy3kibjPHtSVZDaaxz4oakZBl
2I/IhwrwcNJuTs+MQibtrcVtiD2GmTHh/SEp4D2SoRWdLKfzJHSQNW1ZmVQFxbE+LkVp+2mS+sa6
KBTSijZBoAM9Z9alrHjxk793cDl0cnzELgLa6P9L8XNM8DdhemndhPO0HdHrYsdTiaOtTurIvEvO
RzTYCO6EL3pO0bzra+QU/GVRqzxHByPBENsNKLV2uP6gMrhiB6YYcU0K1h2oOeDnLIRG7RSthzGH
KYO5JttZChmMH1v7Hqj/LogJj6ZmF7gNRvOROQpWZLMYttDi2j5nV0ZUJBhxXbL88xIR5l3PBoQL
gNfeq4OPoxZRXEJW80YOO+ZTcWQjK6Hln7s91Uqyu+1E89HLvnYASwcC/QWBCemSVayPV25sDwW4
hbwjFjBibEkXYK8gcgAB4HYNoto7RnjS/8lSft1npogGpNnsRIBelZ1tln0ggCrKygEw9O9WxV5c
lrBPWBfUFbpOi7If2X1F+eOAfH3A93msYGBh8REgK77gZpJk0zvFC6+08uYXvn5eJ8Va2anzf4Qd
YWfHNnaR4y+podGgy/PWF2x34RfaX7krJEg1qekSyrxApyEc3Zj0KI/VHY3I/3aTNJR4+IcNYjvl
xq+fB0hNK7zkoMILLNEb+9QXCa+ZDhCEt0CPgz0iPa4eVkc51aD3m1cs8vbTuuHXMaksITVin+/W
0iR/79KLeHbng5Ytey07TYiYyNduPA8wTaSfk1QF6X5eNWZxevSYG5Yd1Z3qe+c691vMtVjGFY9M
ixL2q7cr4hHbyXyRWFJNKInPrNjn7vLkrTQP58mG6qcnXHNho8SWbC8grSc7ogDmzjBvY0pWyx3G
lKYpwxApAt8IXDScSYN1hJAZ8PXZrtztHpDxxNUpoDsBXryKb/7bVEfGvhXIZ9+WEKLeuqIUKcZN
m9fFQ+kUNZWqLZKnr7+JFBaE3xux0a8XPpqOIsb9GpEQnDRMlyTNFbNqlvAJc8u8XLiVlh+1DVoU
vWpExa6ZJ1DrwZXjFTMS0ysBI8y0YVCCmVrpRon7MZfpuFUkvHzNhT09uEA6YfwX261HaAJitLRU
5pFqhs8WwPdOzXF2uDO+HSCOGwQTFiwG52tLqx59rB3Z3/JaI6j9vYBIwTG5XKn1woT60/nNjC0v
vu/Yvk5MTpuLEBFMIb8ppcbBjAxin9OLsylRqNPd9gqk8K33TnGUsgUFYTDVc+fPqKtfixpK8f1W
cwP8CGh3ct++HKM1BxsWklCRWhNhV0w8Yv3/yhw91AOqa83xhxd3q4Plg2pDRmW24XfMzCkjXLE1
QE74WVPFcJp9f1EptwzBpKljVaA2MuDZFQeZZQ7VkTyf6oomINYWRJA6zB0wwg9tKUlhb1MKCrFQ
5I2h0u9ZX8dJKS+IoUMwABBx4FbthatPIkEDoHez/L/WtazdL1jHRUyYGtXCf7LAVnuoha5tM+8z
gx/9pfqiAd323Jj0RWH8cQkgt8s0R0fuZ6MJQcypf+E3iPwBMr8ArUdqXRQh/5Yv3YmWtPcDFAuy
uNPn8ZlAQqVdGDkNl7OYZl9KDc99tP9p8ULVpf62Bv+jHh2T8rQIaX7cvlXjKL5SyjLcKGR1OOB6
FqQv0yh0uDYj6imBFE3j6FDPobUS6mI9OAn0ig3pESVfGAcVTneua02jtV4v+NMJsh0BCPk7a3dn
uLVb7UO6iJTDZ8BWyaY2MWqInldkHW/xUOfK3sBjBym0ws4/bmaL1rYNbDib8rhDzqfBFNrhesTS
Sh/gbstgeZeySHy1XvdsGkEyvQoWU42jPPDF6oARRx/n9dlxc1juy37if6uEUPZYIPLZwecTSz7S
WDoTfubhQIWRXB3ytI6/pet7YNUbLmEgIuXkN2CNKR5JsWbcWCE1Ptt/y03BVNkhcuJ0QSOUhmXL
PRokCb2z10dWKXXiFHxrBfNKcGIeA4sxnUL+zYxmIOjs9hoS54VFITKT6yB0F8tVnDAwBADYjywU
dlxMV4z8ygF3IEAGQAouthgtlqmZqhx8Q3vIBbqxDsZwx8oeKtlKGY0qMSC7bbBlHFjB5A/Fd3SN
mx0oZylujMMI2erSaYaSGqlHcrzr40EGqTFdsCrbR1BY3Bk3YHOAnF1B69TZ+OfEo8rUhaW6CtaL
FSdcvQlsyEti+HBqM/XpL6p4iqIKZRmBW0hz71kBJZVI1N6he6PbA2rbCz0XEZqeXCGcjZ9DROe3
f5dBIbMUdKkhagwoikr64DsdgzOoALIHYKVQX1caz//7MbDsyUAVMt1oPuU8cjn+mWoy0QuA49Ml
4f1wwhHLhOpDdbBNCMR1doUnF4LfIe0hYczGdnBvCi5+KYGnXnnBNDMbiHNiOtIFq42Xw77h9B3r
O2pBQ8Ja4H5EjKYu9nvgrA0almTV8PgugNpu/Z3m1Dhg8komF3mIcF+9ovUS0EeqMN6vMj0a6D3G
5SedejPDpNTisjWyz7aULRhGZX6pcF0KeCDC2eDAlfJhaQcUD67WUP75z+u+pu5MMVeRv9h5VkkA
lWWrHg4A8Toiscq2cvygetiOlFJpZP2Q1fzIj5CwhE9YAdi7uclcHOlXSPIMiE6TkfoHzb5f5PvQ
JIatdxeEAS7AGYbG7ug0yMyo2X142KJYg1cRn9JrNyL3vv19xdia2DNLefjFhn88bcGWjNFV+rPv
BOuHs7i1l83O9uIkf+fSGybxvx1iM6AutM+P0hs6fI9a7ffapkjh4ko2DFwycWrnAWCUg5Pydw/N
qekth1Rh/6V2rfjZKOfPjwOb4cQoMFNiixQpTN5P3yFJBVIGp9yNV4qpCuIN+0IOjrbG/bQZvcRf
tl0WN8nAJ8gsW4eVLHzIgecuLl64fD/KW4vGeJy6cnbVWQCyOjHhshABgFObHUHLUUYAE7rUOJfh
unojTJJjtZnjUp5oYmxhjXmbQ4qkniyETgSHYuOQdL/qBve8DW4QgUMeqhy2luFigdtJ4ZPfr4ES
tSfxx+D9PF/xrMC2EcOCgUn3ClMynFuMcr5A1QDgECI+oQlw54ADlrALNkJnsRchl4/6D/aU9TKF
eKS9CEDnDEgho6eA+7izPP0EOJ/2jYDrNNKI1TG1k9aJSoq7mainXBlGkS2lY/XVMVNsyKFI7//T
kiDPnMjJWlvBovV+LbYS3HrtOPF/Mbym4rPUEO3U9YMymAJEnDpN6S0bYW/7oYZ9KR80rR+mNBtW
7rTPBe5awwEb/ZU4xg/toEe86BoOa1TxQVMmt/bMHkRTWUO77UoEX/NnBL8lThhlSUDPqc1eRI7j
hCNQUODLXMq5k/Kh2wg3Doj5AlZYkq+H3sL6O4c/d1nJm6AHZYGhi8F+5/hSkcL0P+/aH5G52Va2
svizBIQiqqHBYdp8TngFAeGh0UipsOZL0qFpOsiv5zvpBTEGLN+DSLV27QsdCVreKovYZII7zJUS
uikSdRNT42N2PyPZnGdjG3Y02vvEWomoC5hGHIrUSH42bkpYdwFBWyS9+ZA6NCGyCJDgjiFHWF8r
JOUSLYz6/9aRnH6ILuby10MH4jLsHyhrg1rZltnanNyN5ANYG2ROVhlzriYOKz4DPlVzM+EdENW5
DmXs+jiepCSYbj44YAuLcdt8A9xt648nNfy7CAlOldtUVHznhhuUYU40MdZfen8kI32L141KDNEC
vT7qY0C9n6xTuv70M2jYOaIYgDVyWpBTAvRql+I0iYh2aZjgHqeWs8a3ljOIarEMA3eLZo/yTnXn
YXkQBJKE3e4wAdpiUz3TeL0Oa6j9BCHALv8UZFV42kSyFGU/Hg6kJOEJs1CD1fTF9aZmhDqjYSL7
PcD2sszCzPrZHc+aiplWfc1+UpdD1uIls2jNmB0W+pN7SR3H0+iv8zgajdmW4HhzFEQCq2hksGF4
WrxCD8eOuO7cD2Tzf46GQrGTXIXIMjxqU4CedKql2aoby9KKVwB7yqxqINIg1ZzHe48mxdZ3Y9Wj
/0o0XYAloBYXM48O0w4drbyXOi564QmFq9Tyl9THLcp0tqjZHSqqw1cTSeVsejV75EdSyikTyM97
oG/U6pgVJIQb3LpaSeVSrv9XDdcNVfWb3yOBM4euE8ReoWOEoSU6g8gyTkiV4iSbWgOIIha+7iN6
4l3qFQKshOOW6HvlIQZa3GJE6ukwKS9aRqiIvMiAUKPVpNsCm1ME7UvJ0ZNB+AyziAqCQFgEkG32
/+3oSkl2PTge6STcy5jl4TEMN/JI3LPSQWboncldUQcumD8tWXHudphhPvFBjPUu3LfR3H8z2FYa
M9asZC2GsX/Ea69CqHF/Y5wvdNMLoi+IheaesRM9fdjvoJEfFShJlKMTAvzSdkxvl33RlGqQ4GWX
r+fKjQtzm6/TxhoNGL/mz2CkAFBhgrvIWu7q0zbymOKl9XlAFWAp+x53u9NQrP5mJUNiq/Clh1n2
SPu9r6EPYdcTYVzbhjgdoM0y7f8UNtXjWOcU8tVem7nvprMbUzIto+90EQc5W2PubbtV0YqqiA9Q
xt6KYFzH8W+0deYInGJJKOnMToW4p3nB6rI4lftg/7PkFTG2UJtvnPTVOzi7MyklKPu5WVYDoZvL
uy3M/g2/ACl2WES6IqZY1WST3feG3Ss+hg3Je8JMtbvYVicBeiXfwhAz0gYtp1lyhXkdWv2edek/
tXXE7IVdRlTAHRIVfVWhn9u5g7ee2YJajlHa9SomU547db5ZCeoA9oD6xHIqo3cBlVglYogMXnXK
+HF1VyclLhDSfIodvwAT4kBkrGm1sba8otsKSuBEngc/dDSSDstQ1HtrxKeWoKpNfLB6zwhgMh1Z
SDMD78uFKHpQW4V+fOpd71MIFen2u9b0FDnhRp6HYStmT8BT2NJ4NKFN5W7LOeAbRNr1OK4yRadh
l90/2xAf9PdePCfqgoncCAwulZuGpHqmzuc+QxmF/jZVt3z+zIGiWspO0nO2gbEmh1DrTeBPaaOx
WZQbu7TqvrCSmVBU7s/Aff0yWb+6aQ0P6GgDEBMc+QGWTDvxShOyY4MQQRNkplqZeEu4n4HpevsX
3xeFF2870kEIjiXejwj+47idwBTzMMQL2SEmMp8NB7Je+sM2pVK9xOWVU7MyzISy74dMFjCS4yas
6Se6BGb6HsrPs2PsV1fj2o+q9l131FHuritSEBDpKCLSFpqKLuRJi1CdT/CG+uDpKxXMvp2Rd4Ks
nvr643eo00pWhdO3/vhwLSJJzHx3xepdAiu69R8VdfSZTK2z/2P+wYE6QLN4X/PxC4Co1hZsYZiM
vO7zk4RqSYBwv+/Z+muvPW7w/7OqdrCL2diTUzvJq6PDQtxr1eExVHR3P2RbBk47lM3kjtuR6lkS
bJeV5IHw4s3yWe8yRC8YhbNkFrJftPtF20LseaSV8TeVdcWGksrCntiibIfX5ZxS9UVH0mG4KNPS
komE/zCWjgnAldYKkjLRu1nZf+7hSebqmTVRhhIlNZEgNwrMFRZ+pDVESoJSwpK8/49m6bZW7q+L
OtcfAaskr0mjSFG2ljC7IXNBiBMlytJDYIvICCzfCrovF/bx6RAZbQpW2vE3ZOlYtnZdSOhnJagk
U6o/rOzRyHkOJwSLIyAkRdYvaAK/O7u6E75iD617Q5C6SLLU/7Spz8Oh7J2sNFyb9B2R6MWi+hcG
Saz8LFJ04s+NKA5j/sub75d+zzLvruglhZNc7sVzkUYtIkjREZaZng0rRZBiavfh5MR8HZvgwdMd
UdGRTZXA7hUbkIFnGn2mgWCVPYwZoQa/q5H1B95Y5ShhwQkQfZZjk02gaKznbg42VrrDTzR89Rql
qHnn+9paI6tJJFXAdUBHYSCTw1FViIP+zJQnhiN9anldw6aJw2Unix9oW94fabXM3F6zWibtgN2B
/Po5eCyRnRAIRSOvmgMu2fRmbY3h3Sl+7Rd1ilTpr/W7U4NZvq2a0jY7UnG+jxUXCY+knbDrDx/Y
ymUSSwiOymalTlgp1ZpLMo/MJNXvmXKbgxpFDMzA+oCNlZanM51PDD5MzACacsxjwJWfQCSpaxee
fD7OOoa1giyiyTFKytO1Rbm5D0ANVdWOzS98sIIhMaCtT5gjBZBrBCk7vkdGwJBiMLae9vCKZhA6
uQxTN8+qsbAGHSXS1AQQQTO2a8h4lQZDFYTFr6BoGkpTSWZFqmdH45uYZ1k72bF0LU0aQ8oZLbN/
VBc5zoqCmd2dIebGOxDCMl4xX5v6aGn6KGBM1N/ZRwgfRiQJJF47dGo6SN9unplWXQJ+BsI6+ogz
dyvcQZJ+afaznC6UpAHwcYScJbCmdc4gF1hTrn2TQMtiCYTC0o0kvDI2zFSbNjzPgo5PH12LDC9T
EbhtLv5/kPbJPezYx9Fi47rdJ3K5Homd/YbFyGtPjJdDwZzVzHLh+3n6qbtQ/0gJAbD4u0debiRZ
aFXPjR/7KBEhPiagygLZwKbW4VzLV2FF1w11MGlwDGcdg+tkeeAkYUp3lzq6tmtG2oRCMiSc8Y/A
VAl54Go1HqcHvowh0lOrVLU60y/u+Spn6YOnu1O2T+/Vs04y7z1gtsrWtl0FhIz57DkesIeaOXMp
jdUGkrmp7bZLGNiD7kMSHgtPbH45jikYZCMxomsV63yk9htttpWInekbQhodeXP25BDqdb6zYoZT
nuWlYypb10KIqWX1L05Vt7Kk785ntX/5ZI6VPj8WQJzwtclQ5GPITYy4kCupzCMPgzE8YuyxoB1d
tgmQzoREqbeiYrWF0htp0cCBcTH/pahgEmFGvQuqTWAA6F0VcjADUM76yrod3hVKmA4BaXUj2tYt
1C/iZ6Kc3K5DIUTG5WZy3BCN6Ny+u9h+ncxLTBazLQgtMTMTpoWZ5e4Zl8tvuemJLpQmn1bgliC3
IWwMIESYfEcGZy8negfe35zlB0cGPPRpLiq1nlXP5VV7h4rjVdhe6HbLIDYQa79c2FEnsE8G2ocD
oeHzdF+Qt223n3SPYL8c8+SbLTOGNzVbHroAPTCx9CG+952rMLhRZGaqYe0YK+BN4yOCvMphEsgt
6bnwpD4Vw+S1G5nfpvjvoMZ0ujzZkDv01tU8Yt0sa5nwLr1zx/1maeNWqAtuEeqa46A16R6wNYrJ
nrGc0VGvGdtwUXAWufSfTDA85vYRSj+WZnECKr+XFP60//v0ujs9+n+jp2tzv2vy8ddiunW4bGm1
L5C7G/sxkT/2CCnbmNqSkqZGvb2afu4gzaJ/sEk2qUxIQua9d24lYRsFRU93FOwz+XLWJHyQFmcY
1SDZiQ0L96ECQGxJML88uTY3iGe0JUe/VUebmFtANQG0XYdXjMiITZj2UqITgyYHfMHFp5UfudoJ
81g5F+47rpgGhLz3N0mat+4h50BCPzRttezekcNXnCdu1Kmj5HvBzdvXe8K1LbeGeGDPmAbqElG7
e+gmJDs3fdqXjfd0aFWonKqworO27FPEa2S33RBTOEbYBjGwWAUPboOdGve94MNc9HyrzrKgNOuo
4TMWM30rDCtfEo7dpwJkLRPU1w2x/C04/5xzKqCn6k8o6pCct2jZZ9Dts+X7TbanlcvhNpzqw8DB
1WzjY73XwuKPnX+qTFniClYz8tUGttfmjxAqlzOYh8grotzXUkvTzvuzU9ufoJS59XYJy31ku4WX
wyz56wvVipXbe4lWYeTGROW9EhE4ANed30WNkwYnrlMtAmaSsKu46mvAgKXMNaGT4BGkW2uQmxhn
n3FRxE9tfwvf5P/ZNJSsnL00W7SnZdvZ2T49ik0BIzvkeVZ0RztyKrbqzR0m0ugKPvQIvICrei9E
QUShVkNfmIxcoeEVOqoC1oD5Zs+KLNfmCrREZUAabVnlqjJOALaQhGhNoTq/KLGpX0cl+hnSxIg8
n/KAxWB9fJH/iKzAR4/mexYiqC+GD9CyiHdH1oYveBYrcl2gniP8joAwZIJeX6z39v58ZCqrE2P6
Ut9EvO/GAE/lS+cVdT8AwgGlwTyFmGyw+cHeZFINqaFrDP4ODqANjpYxQULjTOcfOJfd9xd47d9o
7UPb6yBwpE9SnBCsWjP1wx5Vu4dgyN4M2oz+feJyapiEIavFWFeNX0aDWouWvDbQ+H+ypnaSAKuW
TyR2tTzk/YtimF4H/4hjueZ/gw9caNHscYbL8nVilJ49xSql29xLiDruToorpaC/i7L7p963XhqP
q2GsHim9OmJKk/JxduuNRQNx/R5tmt6jXyrTAl2N86hnqm5oKa2JRWDOAXjfrC41LDjggkI0uHYs
/cCrafHKPjlDR1SOuFeStefbxyPijl+ktgk9pgKtWlapWk+TDjrGKcrNeWLA7ELEDyBzvXgsYrHt
DqOeaD1EUJQOPBI7yVdsRVrYH9xN/SDGAcQB/3qNetse4i//pLHZNPUiA9zLExM4flgvbK49AIRY
om4J6+hAZDdgWkYnJae+FwcL0S22oEpKrugywLELs+XLINmdoHDajeKIovPx48DG+0zwONgoKqrR
C9av4hambb6xJXbuuv/6xmVR3duC/XQxE6BoWFiJt0ClDCVwPX8BoCdWDi2Wz84X0MA0mUkDNckY
UN6VvmNNIizn5l+WZ7nhDPkPLOtrXdACSHn4h4aG1tQHTJ3YhhXLkTR7wOQfLvpvO1NIuPCrNtWa
ZslPhgM30jvpwWQjCk/G61qQR/EUvcpphTnMrj2FaiU/LEcLWkf9reE020bNlNCFxBk2hrUdxDit
J+oWVBre6cKQUAWQa733XxP4fQivJRoje0nTKKqpRscZA77TJ2MNEykZuhgdppY10RNv+DwF2Z8s
iEBWnX1IBUIi0KmwU/oXQTsJNbw2nbY41KlEovVuNDjoJzep94OC5CwmV7AleCxvKKJ63rUpYCHc
+4soHe7Ib31am45Uv5YCVVljEBabtvJR8ZMCp9HLN8zDxfJiAWaSueUKsG9PSF9O6M7DYAHxBD+G
MCTC94a8pNExVuQvvmYmPpQNbKucRhJ7vCfZ1Qlbw+UKT9m+GNp/9vKPNyIBDaCg/0WbvdgT+X7y
oTH/iHQDo5ZDITNb8Cp8dPDULhT+aq/DIAO0oXYToBAZ6AgF+hIxdCZxZE0tZv5kpMeT5glUp1k8
U+ZcPtuYxY6z/z4acEgbb1cZEeTTAQdkltvvM67DMDFVk73/tKBgvtxbuT6vAYF8WpkeGv8yB3MJ
daateLEnSy4xfM26vs7VGUqf04QbIT8naUPLdDOHKTnN8zqyddWYMVg/96vm13mq1WoPSvUuFPJ4
Ang+EJlbVyimuK12FfuXDFAV29sq3L6ofFfflCux6TJDL0j6GOVdCyG53JQhiawA1lOrTt/rHihw
365YwFRs720FOc+CeKITQ3XGv2jTz8nGQW0415Hcqyjka2nZWtWA74KubgV558gqOrfBohmlibCG
oQBddLOS+hV7ClhImbJP3IgSHp4o0YcX1zZL0l5xyK3XnGp2bx/bO0kSKyrMYcVqjzCw3aMOHqCs
WR7YV9z2ZijhdTSf0Vo+MNCsPAsxag8QRs/LgIu2g0YWvGzH5aIDqU6Uk3amy/k1P0z3/UoiLGUv
BgpvKICWQqiW5M8qxCgmDRJzc+iJsf/OibMYSgYnqygIIaf0odZL66v9jmPqZ18ZqPc3EtpACUde
9neEkQ8qhKNF3+7BW3R4qJ9Q+2gW66dVuIRol5i2SwWm8BWh7RfLBDE2OEraJllF6laIwtPUYh+y
5G1KVer4RqFNrCqnWff6ylY4YBeCkBq+MNkMmX+foraJyYDmI+fjfMhXPXBGyJwZOLINaohBMR+Y
5Hw2Er2ivmwbxEy88hdhhCK5f7d/QNf2sA88A7JzbAa+b/S1BQZ6ZmTBgWlfkyy+4Evmm63/hpli
ed2XTFdGfTagHucKb9AHsxdfAkSFlNWnUhiEoj50AE4VsaoDpRU/sFXru0c8J5+mOIXm+tO7a7Pr
N5E6Gs61ORznLVMlA8z2mRXXoYzEAy+1W8jbYBo4tTBd29J0Pvgu1aLAjcgLH2ZLGXCRDVERQtYh
vPbi9pLRu6hBLEYeYsBEKHy29koK1Gi9dalOm+QPALG3qoiLGgtRoUimPLuz1oV14ad+SRyltDTL
NURcDXhBuxPpHGZMWSTdEA+YNy7rQdnaVYBhwqs6aCVPaaDVV2ydqeYBLuy558o5xIKQEBXlo6Ag
Oh9SlxIctJRo7Pt5MpDGb8ns7Qa/UKrWVM5aXEqy/BGS8IIiovA3Mc1R6iivxJub3w1Vo0eIswNq
X3jw9DFD4VDnngO/2SWvlmloh0wSZmBDFc5oQLtSsXU2FSBkp4WVLRofRT9oyea8lTKdKgBEyx3d
ja6BO757EEde/WgWg8U72RwYXiU/ABZiQ1JTQt1ZaEz+60v8JyBNElMPv0rZWuLQwby6yRc/UHbO
+pb1vSCEhLdmi3SMkOEjimM2HHSrNaL5wlOe17yhS2XLJX6E3MOdCBaIPOOiajc+TeGA2LefFMr0
DVURLUXYjQP5Cx2zQBSQ+LZIwyj/e1bcmrEbfob8CoX7kdd/pVQfM+HRUbLNsgeFF8aRE7fE2wgM
zPDrYykV7Mc709f6aFJFZB/u116Q1En+C2r3ZLjLt0LWYaJDOYBIE66+sIjhuiKC7p2zl5zAwJIr
Nc91NI7MGRDbvejzrrGEFhYA/U1rPrhf1iIq+e0Cw+wavxRVMnvIQBQFduLAlTOnYnjmL53hjlAG
wlHfkhHeZYn/uva33PELiipUI5Z2W+kFZjHpya52Jo4R87e25q3a+/RKaGhRVHOU0MAYxNc/X9L5
MYVGppHBsH2IrZLY8iDr5UdvoHGt1uUHzBELS+6GW6CNT1qEuM39CzoZlEwDDbIiU2qmoDlDVKC+
i3XrJnRlobeUgHWhA+qJJA9LNf7mPPcVKDhyU3BxwMshdKbmf9V13yglLqjir5S+if/0XDm5nOKJ
CYHeFhaGkZPQBT/9Clrj+XyI5tr7hf9+orQ365dyA8ue7PB0o/qr+tBg8voyDts9M6eQUE9risrg
HMVLIDVxDPE/ynXfNzANqkby0bEY3fis84YeINCnNVrrZueGYZQ093eEFbJUOi5XkS2y70Savxaf
JOOOzbNjelNBtFrvOzSiy7YmPtVO8ZjLO2FSX/mTW73Ga9OSu/yWSivGLY1nYKau4C2Bx7AG79Ml
4wzM/iD3YrNsColAxnoo0vHJ4HFZPtWKU3ggLKRL62BhyY0jbgv743pc23qZomOfBYYul0tQ8G7l
rTIt1A/X9Ookhs8p0HKoF7pkaMa8KqC+F3VPefcZtEPYMLIDKVAqOS+XiYPHb39CaiMe2H+6+bqs
eYWqaOR5SCPrvOKhfZki4Zb6D4w5cslg+KejKkuTfoT0v2SrZWWgYBq4klJFfV5SUKOFtIiRhTLb
GYM3YQta3gCWHFoD9Eg7j1aTZzC5ycZ0yugo+4eHZb75xx5MumqWC0dtvAptjWMcsJ7dRrpJ4U2G
lfSvZxAAQnoHhKGnvUQ4z6f/3TyeMVql2L86NT1Y6sfKrn4wTswcrRVKw3iFtnW+JKmmhVY4HbJ4
KjwlXsMga97SkFxoTKFsD1dlvO5Efa/nitF6aFDvrZAtfzh38PWTuqKbXk/gvlPgHxC5FMZO1EFZ
E77AdPa5YbqxBUaORYbCuTzsIWwQCxqPo7Dgb/gEiwYxSIYR61FWJb5rWhGfMPEBj2ld74IzGL2o
msKXNDYX6TtXsKzNYoqZcrtp5yH2t+z7xVHpSJDlrWgHSk5GPZ5KX2IqyyCewLdYZdzNLYwCK3xb
Pt+05lmj3U23ejLm0JQhcZkFycVoEwXhy2twTF79K6oQwIhnm56hvao0IvysmNR9MaiRhSjVLpKT
YEgmx1H7uHqS0pDAmOMhwo+Q4AEb6Od1HZVr7SqE1OKiz/nZJDYancF5k2rrGkHQYvLSktNT+rpn
2zImjvQqq+3MYTGhloCw5FKto1XlXOX00ImTT2j4SVqxou2llKtpqrCXhjJ8Mb4s+Rmqak5lSIdh
/B0kdoUcf5lQczqDHhgm1ngriw71UfubENxO5OvcRF0YQfvvWeTuHoaxltwBGgpwbJQxbEfkWEtk
r6JRxoghRKochLQJl3aKDy5EWjKycQ6JO0rTt28GpCQSusegwnXDTvrhQf4/oxtbK4GwXk8NfJEj
kr88tHZJ6JLguJRT6pWsNMz6fMeapfQaaONwIC7NVHBjZ7iKUq6O1KTguOo6KbkqUibHn64elhqs
eco0uWCu9K6SeOvLy5MN7Tadz2sqR74yUWPpNjUz/fRuigwJl6WaqrEDDMHSv4r1Tf3TxYHxikvC
JXn+NeJ6b9QEZofd2xUlvdimA+XBL1T7DVO/v7Y2nJgGHKdn1UYX+7B4UrGjp+6nsxAHa5hkq3k+
+Ao5eWkuQ0MU+3bQXksCaMPIZN8wcIFwqSD1h3A4Qi/drjfk3GeNNdYL+TbSJgwszetC7mzEWlWa
OOKaCiblqx0kZUdWnEWOOl9zMWb5fF2TG2NIqvb9uYkNbWwNvD4PZfRPqaj/aPotCfA8bdOVNjL8
Gvb6k9gP7z53pg1YudRKqhK5RUgHVlxDfkD2Lpij/c4hbcXtZu1+peupBCI+JLXGz2j6p507sNXQ
gkiql0VlxjA9TUbmPNH+hyMgWDy3PUMJShzm/09phiCnMBxQ0T6O+HgBWAoJDyUWx6DZP1E9sKug
IB+IoJQVzc54v5unxkEYaGF76vdd7hA8bjWOuaUZlwKzW+vefS77cqXeJ1ROk18fFBZY2r0jin8+
zUWw3KE+e9gNuuvXdZV+CAnPSdGVIeNGhAXIYzRYJeWrVAymSnPZ09FO19eRsTiidrcDT+Zw2k9G
IQvd8prQixmqZ5rKjm3q3q+RaTVb4Qz+fTqzJMd1Kv+uKWNm0untEHAxXE1im8vYrcnOM6N8u1QI
In5CaIzyulcz8C6/44vnWdZ+V7VM0R219WLdgGUulfUr1/ItfUDpjQrN0ZRLtq2s0G0IuVZVP+cX
wkZrGbx/UO+R6xJsAFCRjs3cYRE16vR6gH2IwZ6o/5DRPibKwID55HXS7/oRve2o4hvE2T6yJ609
I6TzTNPaL/RtRPMhNBPS9wb7PlP5HEwVX1gBX256Masp7rdahsW44iEyrFMLwO/8YxqpfskYYhZQ
l9s3RAngCkuaCFa8lIzgwkt/RrbL9fuIsZJ/1ptxDUrZEeZMi/vgMHzFszYDI0HSBdTgIesKIhfE
6OHjSePlCK4fiKaWnlCw2gH/PlmAllEL0lFlYnqu1HlBXBAFVPRg2+8Wlg+miXpZ/wW0sdjoj5RP
t0kgjcAJz3R1rK+US/NguJA1csMXjOl+frtGXZBiQ4AUB+4j7krFgdwGlSAOjti5xG73MMk4KP1M
1xEUXKwPK7RV1B+z5+RYoN6fFMHXYHZxfMfI45z8Iai7JktBO5/LYrcEcvPTufhC3WtJ3fOE8937
zl53vVIN0e+n7UTiwW1xz/R+DHofShNkbSmOf8NHCz1TG8QhXBHz+XeaU+scI+BsDLH91facxPFf
xiXUYW/QnOiQCgS5H5Dn1GAirz1a/Cb8coIDf6zkj4Vsozb3e/yEF4BR3Q8xOmKv+CYaz2YhkNUu
rX0vldb4WJuQfOMe3iGOdG7u3F0oneOow/EEuhLALxVOKlKrvFmheHoFLXB2dUdo/6ZGLozTw68m
0CO2wT+MGngxPFSLWYkyi72F33aFoHw8MatwN/cVD2Hil8LVzvZUh6kMDSzmo+szNj6T18RsfOs4
W9Q3BiGx5uixzcG5Ok1MIYbBX0ppoBLVsW9bQVYvrSfepf8qFBBzPjGkE5JL/lk/nUshRYXM06Yq
0v0uXfEZmbllsMkyydUs4RhEGJ0UBvg5COPpqkeNbCaJ4YCOj3xNPAA4ixb4QGmSXgu1Z7pYWmfX
8Np30nkDdgqc4SwhVfiLaezdnq99CXz9dlylHqDTw6kBbBh/9KYSxDxVnKo7X/gqLrfvJrstfIGl
OeFK4aS8qw60Ml2KJ0Sg4zYoc1gfJM+iRZykfXEVubKtProKzsxmrSlLsV4wUvnwaKCVrQLFoh+Y
PZQytAqcLc4tH1jYsZ2DLZ+mVpMbA5SO5TaKYhIHaTMakm6guVvIApsRnCxzvTV7EV1k4Hg+MK4U
6Jbx432ytpg0q/rtUizHZPPdXsd1PuIt9BBI1meIeoAMFkv8R/Xmd9ZJnbO501UYLeQtUh1oEeoF
az9RnP5moD0aCWMsVze8qfNSiCUH5ujpFzhdXBnNZZL1dRuH+Z8m6plKmeJcfg4NtCdd++H25QT/
tc/Wr6CVvRXJPJMpXJWXsYi35PUtsjLz1Luw5yYneoVYnwSDzEzL1CUDITP+K8M2todz7qtjEtOJ
6N8exALPHc35hKljU4iEb5Zby9VTBa+FuFfkIhvGXrfPS5ksx3bDD/gDqZcRmVy9JTwlq5h+n2wY
9BlyScDUJtyXPiviq4U79RVzWdYaI+rK7X7DkoYOOC1RA8a+lLPEx+KNVru9Fvh0YdtWKEt5YN5N
iB+tsUawPJBm3lc3b3D5oX9rN5qdliRFqqigQUCrWpnE3Wu1Q4yP6EkefE5NAk7tY8a5osvxJ9EI
P0O2xV+LX9ZZInyY2vuaKz2RYBr6os7vUvLCcsTzDsLxiYF97Az6YJo9upoS2DJjfG0k6xPWI7cP
GwJFmI+MhigjUD9KGDBXUkTyvPpMwBd5iHkdEmBK/ouGPnpVH9K/TP35XJZCv1qC50xxccOL88cu
K7k8+g8itV88WyG6C/dcQQkcbyzTrKr1bPacIHpCkAskTSsNj7h4VnxgTYQyYYiXq9xWNS/yNloS
Vymu1oIzUMpjIyfM7xDvK5kAu4sQAeN3AzumADcZVa6+1pzOn54spQToxAeuvzGHIU2PQzn3vpBt
yJCMgfC6trxYa05v/zhfqssGa0zpLxc/odl35i9ifS/qb9+fH397m7PdzoNvc5HnTbiyEKGkQWgk
LVY7AC9vkzcP2aAHwFPTd47MGmTfKpokT235j390mJJOcgjbwie9p3PZAIWJkVOMOw+7uciYWRfd
oJxeUV2gUe1dP1Oh5TdbP5FuhC/4SSQufBbFz+AIARMBvfB8PnjUWIujQbz7aBh5Fp4g5ncL/QNe
1KRELAklmAEeKp7C6r4h/kLXFazLXaFFXWZMAhd6Z8BW0mO6JupVjkg+E581sdgEqdWa5pxlYNxK
uUsUpYOxx1w4j4fOHaoKTS31846FW9xp0laPYy8C3/6AO77EW679HaF5XBq4bwAp7tDCisbR8ohZ
KCUnhCjL21CuD5se53nTAAZ2K0l4xE8jDNwCtsjlTSo+I5yolbp8q15IBWqohSgakZlGYiL95k3U
GuXRndXszMcf689laVTIdbrB74Srpzt1w/pb8a7VV80egzSHZqIjIeP13r1pxhx2qLzu+jZPWPin
n3aXQVaieuwb16G0H4q/kznYZzQMb0dnnHfIWPjwk38Pbj4kVPD7mYRF8Hupt5eFrEViM3Nf9geb
qfECM58Y+gM9/GqWfUeqlOQR9nld2HgVEZuJsfwbuMpK344aYhuxum+P4By03DTDdVk4s4gjUEPl
bZ8FyNKYn99mgcUo2ZhcPEIp0nH/i9kZ6M37vWY2G9/Ry/hBjdwbDG1y2K3EQ9hVJy6b5QGqG0DC
l2XiPp0v1Dszvhb3QEzvnFBCDUXSgdbPKBWReCB345cdEFBFE+yfHe4ELKpYRQZsCcQ8Jlg4xKfu
3umpWK8M5ZKSsRj8LhDDXpfB5FfAVIALypgFdRUkTyYXID78EuRXhppsn0uUvjg4HBV56CYRhygx
CegTZmWDS84J1LZlZfZbNNUe2b+unuEE5sJ902GFFgMDWJrou67ST95KlKAUwUcoaSzkLxhDqJQg
gZqVpTo/5VkXO/8gcViOBghwwF57TDGb0bKIK6e60D7y7vmEijoYAyYSjgUZCwGXSBoM55GOe7oR
YnFQw5kIYc5d7L68qLmR9NNJSKVtTlQFpJ2t4prqX6hYeFx/IDLayriEPMUPFMcJ27Ih07hxCLT6
1/fEFo3HVbB5+sKHAneQgS3C716VfeINMcG4l3JnkFN9EwA/E1ScJ68Q+bieaxnRc7GzY7Pb7Dcg
lNhfPa06AJQ/0reDZkkDa/xhKuhcgeyQeiICTW91bmF3T07NAFyXtdSXQxoXR7tGAGBE2gztXy0b
xtL2ADolkIsEdZcC72cEHcqmOUnl+09L0pkPfQVSBz9ZnArYXUTr1lOfC+pTkLa7RKVi+zWf0nS1
7kGSu1WHYt8za1e+5aYSkwB9Dw+3zigSq/YhG3K0f91CXWQ3tO9RySOzA/Kug3qo8gw7hwgesOkY
Yljg1bVNIOCWOk5JGzddlBfyGlGGAXyUoVtJG7o+m87Rd+aqX0JLeFywxDejD7KmGvz+byDRiVjg
I2Uhexo3tr5QX5HaUPKiz2NLAVeyt75thvG/gbASqlXuW4Ld/GAGMCXVqQcmM5IOF9qNdHoCZkSK
r4tGB1ck/MV8gOTsXIzbtXnnMP/fL0kz+2UNi8SILvlHdn1b9HzL2ho35g97QDO6FWQW9FDuasMo
C3iFtlZTzIQa/ykfpoqRa4Z0TTWPb9rADrqySvdiKrSbFmDyCLpjl1E3TOHhXbE8Dz4jNwUes5vF
kiDJWqfnqGOrvORiQ9pUVxUSqlPcINB88LP0AKeqGGTPQQsxeBVamI0fPZhz9mqIHJmLhWBXTPZG
kUlXtCAd/eT7Llw4DUmwgg+EPbeE7sdKUg/JLZDjtvEHDDMSWxtA4Q2eBFpp5bSdAdxKSER1ZS6a
kxwSF5J2CnibVbU5v47ZoSljnbtNXcKRecLvPdi+1iwihphDTCvtJQeSJWv5XNITYTRo9kOhtuFU
hU2aKa/4bCicu6xlJ+q8Qwv0qtXNapLN2z3N5kiB0ag6NKytYgYdbqc3CwAhNESoS0SANJgy5Ou1
jaC2JQLFEM205fPiBBcr0gBHkuyixRnY1LwH4kWYygL4MWmt8FKAFgJ/G5ZtwPVpY9b44RyY4iYx
AjiWEqAnmaj0mVff1iQr/5xZyQipYM8L5Y+ZLmViBLaqBwIuTO5isH38opjvixHl1qyWXirOpP/+
QSl2kjrf3abioV4NIfDGBqMZdJR/mBv5umYu/JoNCePpIHla+TBWrq2PQ5f2P5t3oY6j9QNMhP6j
5j3BiyjuEfn9WQyNj5KuauDK9yyjyGKlZVvYf3B9V4D0sA/2tB7VQIJb0YhPyXf7lm072+2CTTpf
5KlTYxtFF89jBLXyv8C3FPlgTKuhL0zx1LlYJp49Q86fr2pOAAv4HVNNZUfxt/Aqxx4H4Oxja56d
nNgd5+g+wD7yz3Cv5lz/Xi4zI0nVNyvXLNjyPfcWGAlOAf8Ly9mycLUmfFv1a6jw3jJmUcEaTUV2
qReTQxDqiVmc7d+3yl/xa7uU2tYxMOnOSk+svEO7GaNpSWxHD9ASM5bkq5A1161w9KWDwjRjbHDu
ee42T7qvYRO4bPTBgdMbacDKIg7O4uN3EhzIIEXEJM/wPA6AR+g3X5liBwWOzJFLqkHLh323ysW0
sTmmwg2zljTEz+WX7AQsqd1Fsqux5M4R2IlxRy0gqE6rtLLKTKMDrtvhW7z8Zvph7NRRVcOCWvGD
XHI5VJxdToz1WIEs2OcdEKV0dOvnQAgPUTXn50ucVXNR5qsU4+56IfyEyHZFk3Knv+yDu8Q9udbh
J7y04SWZyS595mTAmKfaBqUBMPsrWcaloZp6XjZN6gkDtaymoJvSyeHjAaxfqzOiIjPVFcH2kXYS
rotUOjGF4aWYrIy76Rs46ki5kfbX3MgCypcenAUj2cifMUymlKv8XNj3GKA1Nq66H3idDjA3mGgd
gCEPaOh8YVZSzxBz61MvYN8M8RE269UTh68qZL6RGBjd/1uFG7gV2ck2pRDcAdZDiqcQ1/+UXZT5
r7ZP8LWGJuwcRrpFpBJkQ4m5DwO9Kc6CiqLgx5m97jQEUtCshWHPTvgEpuc2fZ4MZEme1SpiLz5t
KuJfapAB56cXEOYLPKiQ17xerSgMssqEpjD+eNpXGKwjoEd/3YR4fg24+Gm5TY3pjpDqZAwBBNlg
qrWUzxt+dsXaEjgBilwplC6T83BnaL1RhF91gRERwfzjSLzY7gpz/NCvnt+Quk6qo03hv5JVpAMB
dhQWY9nLKqzHAb5VRtInqrMJXIEyDDC5GTte16hwn7eP5luaQi323Ss7PHzG9B+Jbxbv70YSi1ZD
sxX4JR08ZaHyEXuxGdX46JeXzM1h5fie5wO7b9sPipJU/YPwwOxXvw0xmRTJDAz8h3mnbSHZuU4J
FmoxgkFe9NSjK/rh4JFnicaiOK6M4GW9lhVM53dXz+yPtSdCfaA5aRs/i6wvrZlL+xnsNQRCVmvC
u5s1wApepTXge5w3gWc77BNkRO+g3P6RKUNZpDYFcl66xHeMlVmfuEgeqvvSWO5UwcKFoK9IO9wa
Pno1RGy73VoC850bs3KOLR54PqJJ4YoHyir6FqA/HdO8an46BpTpcebc8t7peKCFPQxeGiBt0DnV
0FF1/InWQPbwV54HG4uBxjHKtb0LK4mhGXU/AGGhoPkn94qXL+/jIGTDLhGV+oSL23nia+snoBHX
owdWN+ZIiOXFocVjF5ZYidR8osYCmsTwT1NZfFwFAe6U3qm0fk6CMenywcekrBcpSXM3OCJEfCg/
X97BRQECL/anuqdAYWFYx2GJGF6gUHENjpU06oSK8kxEBTOOmaW/qA4V83PhGEC0uEtFySGrp8qO
QIhvGNWe6GDCnuIdaNLYok11TlzuB3Wi57SSn1TQAfFTG+8m2KDMgCrn78T2Hl3+MKvsyxivzApn
RjWz0l7iUI95Pv1MIDL65Yj0iSbJzEuizyk/8gLOB0mlNX2FR6eGB3abHcbwNQPukC7CN5N8hF7w
KFC9YMLsbbX5THI8nWaOwStNmT3l6+B1BSf5sw/YPnJIUb7GEhZOQnROc9wtg7otaxhjgJrCZBTA
AwzcesP5Bi++WhqmDXEhKJTGlmWlenpMHUCF25lA9MwWSDP5+pueOTG89iZL3S50T+p0f5Sl8tqB
gne+72nAXkVq6ooj9qeD85+NE+14otvmtMfAW7Fl87ZreMjU+z5rKxiLO2tuqSCTOPKSttfghul4
RFTL8M5ZnpxeCuCcoSahWxV6hyUS42Qt5fXVIoVUXktqmIHxzGtghp9vxjwCZkhFVwV02J8kvcsh
cj2BQ8bKYQhvRijTs8JZCO5Gbnj8D/IBBiqLP1BIuGIDy5q0aaE24VvVU7eUxtApBAWrb0uDaoAv
zDGkCWFK3LjrarGorTZplfwpcCRCisZ+g+GixdraBdEdPd2VpjNHGOK4Uq+odQ+VDx/VzuUesMEB
5RFk92il6q3pS1kxpsnoYBhXRvajhduLRibJhsXaOxBNMNXq7r9UUHKZjk7szzAGiIO3WDxxiIbm
UtaQJMPZbR6vU2VAyK6C9ZW19neJA4+3+0pLCx+aFGSJy0+FmvuYT1S+2RMPlzhzkg2g6bcPfx6F
5hzvZc02dwrOCu2/cVSxtQgoHZOowVcPptEejpsLd+fjuFfKj2c2p4AcMHDKoUGLhSu4K+tMed9d
fIVZSh2qMMKlxYRVtSqVzkr2G9uOplAmbZO/UsYA7vYkY0PY/sO0vYiErD1C/I7uQYXhKFkXvovP
MKx+3InGrx9nO6R79ybu5hWkucCXtjeGdEGSHxe8Mx/8KsBtal8XHxTz7L2+/apTViuw4HJGy1SN
z2k3YRasH9MmzA2Okx+45E84Km1z2lXe47w8TtYa1oVJKFJo23dNhkIZu9T6CR3xz+MiCFAKTCXf
HdP8lUxjHEWRmqHREDi0fXpISDfdrVey7tG+DniRc2d3Gf9e4yvuBIrbb91PGlOlSFSKTvOsSJW/
yX3jsg91QabJcQ/FcRw3XKXWJK07lE2nxZoTr340uRbWKmE7C6If74Wv8/Lqg0JyhzIn1D6R0Hg9
gUbIBoQhN1bB4dZaE+noxCROlcLkvGFLSAehL4Z8wWonlXAsFJ6Fj+XF/QSOckyC+Y6dFeaVNPI/
xCyRduCK1awOL6b2YfW4FY65iHq+OemWVmdPvZCnBbmtQtAhH+aROhwQsnJ9bAUXL7eDpEr/5hQr
/cu71pkPTIhCrOjtbp+HcN7xp1UURAv5APmkq2t9Hzy7JBk9/bh2l0NXai7FxIsYUm1feTJ0TxgR
RHTzx16ZUX3ow2VjLyMTU+ehMu3tQOP7G8w/JCuqHWY/c2d6HwjOOSN7ybApw5/yigKlcFHQ942f
rfZ4fqWjy8x5Ij5KgGQX6l2IweoBz2uVix0qtrPfDqHMjb9Go7Y9chtZ8rpPxmE3w9mx2K01uzUE
Q+r0cdVxRqg40XKQQm9TD+QeoKXHrHWDYfxIep2zYA/2ViGMa9kQdVCFr1N1InAf5ta6tJ/MRWQi
ryXSRwbyhh1mIAsPDJELsEr36cjjuGapxwzaelE4Elcgqc/mP531HLYnFkbACQfxTUrH+Q6VvDHz
aQE41OsKXtZsD7VjrFMzRapnEPJN/EN9QnO3RPsIrlpITS9N7QRbhcOlKHyj4EET2jntSXwCvd66
Hq+fB7Y5/bGWpaKQ7V+02FlT2sCNZ70d9zn0RVJ62qfuRtw27NLvh5DmDYJourVDOU6FYEg2u/uD
gRSnspNtexxDzjazc+AEC7GmqFnpMfXyeLv//4WQcfslitNudjbcNvyVytWFJjy1WSySqsDQrIv8
vAOX90t4Qqzo69MP4y4kItpD0vIyNAy2uU1KWjELiQrTxINWLffHi9aPtyMthfve16b0/NDZrX8G
8wSrcvKdNDg3cqEq7x/e9jUjkZ7Ps+Z6FEENWymjZiXzI4BFl8Fl+sRg3hi3dQMHU3h9dqLpRYH7
SJmHh4+1lRlX5BVKhx6eAQJrgK94VG674AuHojTD6B0hnWBieQb/yDEzkM8mIa3vc9qVeJSmRGpP
gwz/OTwI6icwecRozYRh6/Nnop4yYF+eTTn8KuuTggun8KbacOmSjhvjGMPc1CFDf2gufemlmRq4
8upBhloIv+vo9gz99xB5B5WnhcI/i5cFV26hl3d1LLu4z1jH0fvDfUqsAgk1RgzRCPyKbTCCuVrL
g0T7MR3IhhLGQBK9ER3tvOpBWhhGR0DeGuEpJctzAsNPxMtGOGTeB2ec1+QI8kmSOCbelyUpIfTF
A6jI3UvjC+9T0nbL9tTjNc/he5nivwyCNHDDb4yGslaMskG8ZKgL3yIQgmXQ1AjLzf+CA6+jhmsH
NdJ4T9Jp97oE+rZh8oTx7rskfzCvejHjb04q0o9wbTdsmcvIRr+GR0GSd7vkSoKV/ZGt8CeJXu+f
EeP0X1ipF6IctMomEAySTZGurP0ynRmPo7L0Vt6D/Gi9R4GO74ocZwD36CsG+zpz9NwfPL7v/qzI
Xdl2SxOAAsr4shtH81aMGoBnOikyKx50sbdafc5qSlRxih0PY0YEYhjYcd8Df6zEtAFBk1xioJW6
uxmq8gI+1em7qA7s3WwKoTpnPPZNtMuY7O7n1gzFlRNcHoxcZEIQ60WGwMENddvdlBp+ms2lHpS+
0eda9mB2V5iOCGsaOemXOgnwCu2sBOV31PjzXI/igf6IgFCUF4hklywILwlP8FkN5ZPvhiTmXD20
RbvR3PgeuHSbD2DJW0Y+YTPOcZbZGi5PYBgh3PGffbO0/7HQtvYVb72W18tCejQWUYv7qMsU83n4
IEpjfmKWVjDcDm5A2UZMVSRspzgtM2Rgcc0TueMilP7BZjDz82RURNSzWWnVtiU72n/aakVM+CZ6
TqX4G5XB37DUt9F1OWUgZ+Xe/LSvBvhm1Y0+26FqhLZ4H8T6EOdq2ghPKu5G5entRsPJjEY5jn2C
8maBrfW0EctbpWvFZS/cbEAjsqeLJNImWRp42qurn9qyv3jcVoB5xfgNZtekqJk/zgEqiBHWbiG6
77ZpOPGUPyatI7a8ZUm7IcM+vFWwGOmIRa4azX1Ag1Ou2L+zPfjpXU+l+Cv2pCdZ6SCHIS6dwi1J
JzhQqaOnxKnDTPblK3HQcMmPij+aGCkuF93gWSjP6XaM2Zx2twHq96HpA1/QjP/eIoUORbFA+2PW
rDJYF8n3VYkWriKFLMi6UHH4qUWnajGSMa24kTQx35Qs9220MNG4NaqSEvBBhGXj7ZRQCJnlPpNE
84tKPcCqSLrfbwh8DV6afsH2xVSdNQ1cqtuEF8hwDLQxE1lRCCatvIm3MaxXLcLivvPtx2vZr+gh
Tdthj95iz8WvYnZDuXmkG70wa7EgV1x5ZNdTKHhRKo6KNkJyuHt8Us3VuU1tbjKyauhO9c+hEiLj
lJDwNYskSsvPWy0jQp3pAHD+zsqX7niZcjAfV8XDYhIJOkuklEkK4HZxv6qQ3K7vtahvoAm3N18S
m+hIZDrqH8V4/E3G6vQ45gr9tjz4IeMKX0Q/ysgLSK1erudmg88YxBFjQ0igrF4iiPt9vNuow88R
fMiFuBEiLKeo3Xhr2BHwUqrVwxrlpdc1Kyf18faoP2rGlQTn259gLzrX+sPFBRCsRxHoVEQwCmhX
qyG17VqVW6Gp1MSYPd0vwyMpLzAeluJwvkgOe2Qxx1+v1486xggfDtT7Cb3dBFAieS6GNxyses/+
INgr6B58DOoFofGtC1fLzhvSs4EOEvhRqfvL6WNKtyGtoh7HwoJ1y60jat/dOHfXCfRBxi4K6IWh
7AP6FoH92iWENG3cgTCyxanqIC141f4NJLrRfDyF3YpsCBojNSI3HMHUp187MSy6es1RNK28zcKP
/nnMFAdqnPJKkabtfSR1W0SgAxV54cJZeQs+QwoBC96tIsdJRqVuR745XOlTeLkbNtQqCl07QCTY
1VEYq3Pg6Ci/J2KbPENhoz2fuX/eC9Z86/8Lq2RpjWFnLH0MCFKvfYiOMiONlX/OC4/hqrawrns9
xbbzS2QuwQ1vYnTbB2fPujDB4/U/qspqOGtiTuVFmHOVG7VTQQnkSYNr5B9JMlkefQG+xLZeOUK9
2AAsyHaYmfIiSqUBwtQjdlkFCnEk6VnhFABAQqwSdagGpfQc4Y7F5g9jScYhmBKuWwHdudEDIbCQ
ZtaWErKwcPOuSkwk5a3qF2K/hiajYIET8jjT0XRSKkUt8dU41fMGKU/yrlGj7ceMPYYy042X2QtW
FpnSfJ9QDJZnyy9vJPn29adny0NG126UWIxuJkRODW/bs/12vVUDQDyGK/tDwvVOKljpxD/QpXO4
VyS09XTL/pEUA1beHk9gCXOtY8I9IPt/0YWKAKmwoWkpeS1ZlhYAcDhku176FbYBYnYIk+CG/zez
Lckd56w8OCtnmEEucVFmus3871l1+q0Ge4O87zY54r6V4UgyTiaWKkSpWAHjAByozrXWpKNZCEGh
m97n7BSkrYZZC0F4FTb47gVamxk7u8nLHMeHwD93JSwp87ZRYqbOEsu+2zMG3arGgfyt+Z6JNiMa
L/rQh2Epp6aMF3k4wyVB5jBxRrCQgGoeV8sO8AVj/Wtl+fI5sP9iDxilyfhVmPblFx6rn69rXm3m
ws3jgjwRu84T0+DQrrUhVO/AmImuPPv45FWPqHAVQrkY79mvxkUIgGDfbFnN9m+PVHGml+n2WFwd
0P09CCtVtiPpoi0S1HbTU127RauSP1zcfrEWx49iBI5BIfbuESU5K/UOmg6v1/CLgEUOpzPRTf1N
ES3NehH2P7EaFNSzIvYmXV3V+phZ4/aXYmKz3wldCGQthTLQaDnimhmgKgpeQObewfvW2azJdg+h
jBAtESzR6l9HSX6h8G93HPqSbHCwPUCwNJm36ZplWYsoJyB9H+DX9qZ0LL6E8T6iPPqIZr0iWmJa
q/EEVLeIK1NGcGUoLp8pq3GQy6qGG3BEZSaBpQZhawVnPrA4zljCRPwHJcmhPr5zqLAD3HHDrsPu
vl9qXYCsVERGkAuj/W7cc0SxgJoqTI1zsbhfWkFmWUQHZWezcI9iSPsCOnPrCdV7cldsI2h3uIl8
aqhhSDUhJFtEJCUQTaVnav45Rx0NnUY2Ut+cWOPxRNL6cpe/rBjmriL5BcskLugoSvLHhn08RfEw
0w5tjCn4M/cOCbtNNSPC9zuSN+z1RdRPiqQ8Hu9MKVlnldwidio8+JG/NuvPvVhnJ7LzsnLTPegR
kGLUfid6bGKcPjWWqcygigMGrwMUS1rvrnKb6ckCIqRe7nMNLl6C5Sf8HMWhCUZqXS3vc4QCGgGO
L0U7UZJ2Kimq9INtXdIASXPV2de18kQjRL7tugX5sgxicJQU2geOmgHaEPxNfFRsbF+Q6G178Bdl
laZqKqAbpVfM8ULxpkIAmkzxueh7H2LRuEjMbCDdNaVSR7lzy7k0RXx5DNC00t3+Horiib9qWwj7
hLVhN155OVMXAOKlW9jOwVV5P2LFI5nJhjTQU5VBG8HLVIGuBaNCFnUlUki+bVnR2c+W7fHF4tto
urpiZKaWktjy1tr3NPs6q0CUjEtMHI0smkhGIyPIu4/PLdQGOXemqRV5XQuN3xEK8qYQuT0QqRIA
9Ynne/+e4Az2gY4hNO39Dr8w8vRyHMq2t/7oYdyNvyCIIUjFV8plWU+v5dpDaFHNG9Ncl0T0ml5F
XrXwMFrY3D4lnpnyTEiEz4z06jm0fvP+hCZQbu/QN84xOK8ezMVJ6L9IGwTfgQg5qqfS2Yeet+nF
LWO+LFyINTe9Mxvu5GE04rhBkoYsC2It78v7URihX8mKTCYY1n4lsUtkMFkEPCrZH42Z91AW67BA
QS/JHYzhORmcOnwtP3IsJMjW0H4ZVrhxgUUs0YLHOwOmUs9nA3BSl+y0ghnElyf3XmXQ7GIA4NIM
D1MykxN3mjtKnKxznh6kz9WYkRM0g/i5pZ6kguyJFw7mEvMeAbe+bPTgr00K7XlMhMHkWt0nq/3q
7sOvV7siem4mZc+i1Yd9EyqkEBFrJ56uRv4pd0RCh5UdXq1C5aX+nCPVOjp5nKlkq1KxO74WIeSx
1iRwvoyPm/mSljmtmpUYymJhDFhXccQlOD4dSf/Ja6II0JthV5WFocyqPfw2L2l8VLmTL2atiw3D
tTVPiK1mvTNDzKPQH+bitF8V+nuLW9yQGqSMgC+4nIR8Ik3bIL1ISzUBx0nxliNVyo4hJteb7G0l
BMO8unknqzZuoyCjHo6HfGcO1n9JvhBtEkU1VUKaXheAEY4s8iYHM1QyWrWON6TYpKEf0znKozhR
DJAxbafgnBLk4RGb1JNmUJYuL5JZzbEsghAKIKMQrhy2EAAdJ9R/75FObW6laHgh0/Ot4XDth2Hi
ixp6o2g8aKGuQ/bUc5ubozOVw5Ez1wjFmn9rWR+KFy90BhNQUIF5RVKy1zb+hSfgYhJKjsbCueDi
DOHA92IEelR5/Z6vDydmiRp1nT+EZF2ZWJRW5iW0I24Dkp+sTNr48LWg+eY4oEk5MzprUOFt+9m6
cwpjOAZauIwhcdgiVfPBPMthLACTDjuUrjOJlw9v4Q+2xi0ifSCs4nGe+AkFb8kOmM51VvKsXXYp
PkMbds8KB5qHdo7SBDnjy1anmIwGEICC336ruzDqCPNUQ3sPQFF0olGGTB40wZ3zrQ70kjaTUbbV
krUJLSlqtneACBegi10xnqRn8PBQzxQD2ZyTyMZFgvQh1c5v+iNPmUeDBbEND9kmXUbVnbI/IlLA
B3rmbm3Ew6pZYVEiv4Tyvai1P8GN6gb+9jVFqrden+WFYRiBQy1YgFDVFqAT+gpAj52QZzdgVXno
kxVnKV1DN2em4wOmybW4FO2hFrikufinQq4Je0jKM8bbsgEMDoy/WjS5IA2fk3dMYDXJ729t+Dx5
nRWH4BicodlhCrxORn3iv5X87ncI3UeY3aNA1n2vPssPFNt9icCEoXEED5OopiMk546plbpMRURf
OKVzONS2UsFhIEbGnvrQDe8CdruVHtQyCxbP1GGJXNIQmm2PNjQ42PtfsWoPb6BCYtpVhILISBcU
cXhjkehpeNnbi+eI1FeRmfpGFV4l9r7KTxq5L1RwBEQIgOIeV1nAEC6NO6stn/pAlzkrKzA5OWMR
eK3wfdSEJY/kmOMM9Nw+JC4LI57VNe16HuQ49CdPYsO3nSkcbxbYcT5hNXqlxGkg+EbZr0tzrfpo
1wlgMDRAagr50CkGrvbYms1cjnuIDyN4blj+IuKicnUvyNe+XbLJiuqv8yNWMNAZbpGl2r6b2ezu
tH4oje7kHrWUmTBXgtuX7tfQdQdtkQNAouSLtR7ikB7OvIblNmZ4K//QKodrc5TpP1o7TNdTigX6
RHy2g3zW4zdbM0V5hHvUd67cVpSJqnzGUvQWjFx1Az5FR3aFlq0Xwlb3UfHM5ey2RHgxP84ItTf5
Px9AhCeUMRHClBjfvioQpLrH+nqjwReDU2X1jhS2vsGO7w244uCD4ZBltBAvFkwgcuvj2Y5Xx8d3
NBBRhEV97vqMGdANCLd7+hG73Q2axRWrfgQE3/K8cqwTx24OheOIBx4mmd16vZgINZMusL0vyZiw
D4l6gvCoMs647HzAdBuGPW+sgbQ3pOnoUN6ITLiITsh6bfO5PvmK3oER8RBIH+PDO/6ETDisilch
LQK04PWjPbl906GkTt8uO1WTxA8SJEEsl2yWgHgDvmWJVzJ7lXI9kBm4y6MStVWk4LyrUOpHjM4o
yk1U3uN2ItMDXQr3qzfzfoL7c/hGeqhqgrt8wThGFeHvZrPct/G2LzcFwe3EazXQFWQ4mvQuWZN8
9dEJz4D7R6FXpvo6vzEBd6bmTg7aYLF7oOIp5dRIQxsPszv9A9I+jEepM/50+FaQ8YudMr6hm7/L
GCp17/4vaiI3Ewmhljik7kLKTYhXw4aHfYWETwPQv7ik9vIEqULbpAzPdd47hwljjUbukQqskLVr
n94K6PXY3UHWV1AXNVLERTvvQrXJmxzszntGbxUm7n/Q3D7nHmdyQk85sU4Jovu0AeTHa+psmoHM
E0K3+mrqlbewaXF8LDWxQmcXevkdupUI8ajMnDFmeIzQrzKF17xtgpetrKy9/TYgoS9mBpO4lStk
jafvwqnihBakFxcTvfAf4ZRjOyB4/XqlE1Hd1/mgoo0i01eQtHibSgWFIL/WHBu6VeRsqdWocRUq
CNVAJEJktxsCUbCpnVg5c8WnkpdGMTHECGJApq2vcM7XOJD8prueT9BuyrEAekvI3FqPqxhRD9G7
9nSLgUse7S3GnFCGB++0MbQFAcMoWwiVXhqoeVSjBKIjTgO0P3655VKiROAJNxs/3QBeqsxpda1E
q8jlpgIbeyOv/uZcMSD6cfqSx66I0QiWEFDwnXaFRZVm9+e+PbK0D0OuTYB5DyzEaAlGs5o4G/So
9ynYTgKNtYWy68NB17+NfnQrnihm/jJ80gQoUJMB1/7eAkT/0emOwj1Ke0poC9R3o5AtegsfEbxv
KkNEiK+FCtVKuUbRvNalFdOFNlfAEJfOgbdx012V2WkymkJm7PkPfyzHdStu1xMGzQo8HpXI1089
5a5TXG9z5bNCJAf8wbS8mcXDHfUEAEaxXplPvgwrGQgOHy4QQwyS553FWcuvp1lxYPZbAzriiA7V
vi+986eeqTzhs96wdAz8zovUDogATXYMDRX0vIHzAYzyEJJ7d5P8jEHQmeTO4lWHC0UEQSkf9oSt
WmSJIVD4ANKgHqrk2L1MLwGlUao8NvTCHCWZ7cZ5gl6x2v53+I7m+W9fQakfntTNUGLdWoM0/T/1
4Js20kGo6M9hC/wbj6TZBCjebuZp+7vxVQbozEdw3LfgZKp4zkyPjq4Kk3cgwjMdNooczcjfq3Qr
uIX6lr+W5Y6F6uHpwxxeQuv44RtlCF83B2cMSAHm4GwBDL2fYFkzRRGerx1pJJjhVqVp1mf76wWR
eGICUFrFT+gm0PC7k9Fk2mQhKzj6tMV8SSXvotkiZPrmxmjYxvlT69irlFykYSWgQsX/eeeyG9hl
Y6zRsLwR8y4EjUmt7o3tro87LajUQiREch+XI9HkxKCRt3CySTAIpXGxqTZcKKXqSLp7cDHV5HqY
CymIlhS9wdCmHoN3diaJDNTMmniD5HGWPBFJU+tIVXLz/WOwH/rBbAC+MdrJrUzakpajpvcor5Ol
IpChplvDHomcmT1bYMeMPtjSIfyLEomYD03uV2uryBVxmaPNnIA+qxTagtuf6Lc/5j5o9UNRIg4b
fB1wFIpEuzs2bdypGUhhFKea3Y2eGsrEZISHA36QCO0xlTFVzJn4ktamACTSBckGpwcI9ZLo6MIN
tg/uylIAdTI7xJbDrDZhG+4Lj9jE02nmf57zwUtbFz6kOCV9PaKe8gQFGAC/nEBOOtbOlCbDbPAH
EncInqtBBudyWdFTCLpMgQkedf85bP5ZygKnxhfjDSX5ec+pxmY2oKwVya1g9iVZplypP3ToMb1c
MDGy57R7+hkFeiyPdA4EotyCCKHQGs0l4SYlJpnJBpt+PelogOhSbzR7ouGM9s1XTZoutK2r1Q+Z
boGZto0KlIapaTfLSo/GUUBNAi7aNhPshahhxnNbNkdvNZZdIM1ujhImaxihSTyhkC5KkyCFUT80
lyDN7IidwqoPJ6TdrUM0DQx1zDyB1/23rA/W67IhEuCk/JVnN1DPczXSMwB2QhfUCMdZX505Kdcq
U0ekE6poKfBpFfIGUCg4afnBr7K/FHRJVX8HV/SzvbJkqO/TrGoF9/wJ8psrYM7hR0x2JfpkSb9a
4yCsXFBQ4eiSk/DkaBTLU12Vsk6CI+ygd+MrSGyhFCAaYMGyd550Q53VJgPsxtBRlbtWyjkpmj1D
dHzKrKWfcs0++35otP9lMnc5wf218p5hAcH7zBwFcnxlYpOnUb7d2ezGsA1ZvyU3/pnVnKZ1qmX5
J+lDKJbbUZxe5aqF3GvfyId1YREP9n9WdHo1+0nEVf7ALaOeI8tqC1mkdrEibda4nPRRevb9XmzV
x/4QvvYgSHu1qq8ixgbuCMMiXdtMnZQxAs5w0unoss/SflvWZYTVGGljlgyRQ18H9lwj9tkCFonf
KBYjgh9U98nCqWRl2/vu2wRzQtNxSfB0JtQfjd8Fr3vxrZvtPvSTQLOJSapRNlNnK7XvqmgIqa4I
y+J0CwtNsvGDrLim/aLXLDZrUd48eiLqrb3rN00tPz0fcziV5Z6znRRyGyhUf3QIjVz/RqRFsm5z
JuxZ8yCmTj57qkvXpW6cA1LE6GPy99SP1XNtjzAylLcGamdEpYdl//mZHnUM9c41rKXSIZJxx/Lk
LV9vXwHX+Wkp7bFaJS1OneMZHVJIguS0rDhBfj97Vf15bXvMWWgGxSlAnAitPCX1+yDHRButP0Fp
Y8qSYfT/GBbGY9B92QPT4BTFRI1OiVKAqzirLfM9trDpWB47mtX4AgEZVrOWmBtNpNEQf4CDq8eP
koaYpQCWLSKTJfEXb9X+fSkVTzxADkWzBLnsLCoJjg2AmR8nBW21N35IsXD/IwXB8sEP5VKTmBwK
vQBoAz6H+2RISuBrc7UB7H8CLMW7KjKJkQ7zjeJw7Y0szIyNTHfwMa9hNSuNOiAHvxIKAAmSRtSm
5yBh1gtxQjli3g+oq66sLmbcSoWkcvR7Xz7iHWAMoR2TW/frebYLRIIJWcifpssjXF09O7eJ2jyF
l0XIJpT/uJoZQ1oLUzKXUKJKyHJMMjZFkW/z6DjvPFRKmofxX7D9yCk7N6gz6X0+sLBFgKhY6rlm
YHZWIO/wnKfsNapUW/BhOlISJxdDLcgB10k6Q3ZmlqmfQeXRBsh6fqnRG7sDWIG4Kctbw/iTYbws
nXaLRKCcpyGeNZymJ9OIcIt87WOke9nbetnMfQiLv7LBxRAwJlTLEgP2Ge1Aj2H43j4dTEehWayD
s7k5lC9gkb5FFyyR9widf0ecZW4ZlDfkqXQLlTEJ2ebUKZrhFBNvWnzEEY4I9uuVIuwLvsE2Pwf/
9JHtH4OlJFKQ3RFb0MeD9wwX2UjRYkjrT4LceklnH98x1egpW9u9Gzv3nvIiEbsbahdu9yX5lubB
Ywf/ghQiwvOAbj9zUw2M3wC3ax2s2YJcGW/ght6IzyYoiT8F3WiR0Km+lZmzkZihWaM+6DxefJKu
yWHbKRLun9tcaAHqTAJN6lOFziuHjvcoGXBWHZPvfvlZsJpKIhr2iK91PSzBKlYPQdkam3z2qTWs
xIH/6QpM/GOUBP75lz+pPy2vDrKEJ/UEnJwQR1z27OD89DnRST7E5D49+78r5kT4ctKAPstRkQtf
BXl7IqqR0wiJj3t5kP1X4FmKIsoNlhhXkLU05M6/kfYZIBo48Kw1YT9KjJ91jGE/noOWjStpRgd3
1/cRwFAspVA81zMu+zAMc8+lHB2ikrTjblT2ThOJlnmwmWKz49hN8G9zXce/55TjdULD9b2I3DSI
+hUvky4EvQFiqSRYBOpndLrNpd9HRMmc9ePyF8ojtiYDlR81JatAo96soGDGlD0F9HTBRYUVq0Dv
h50Yzc4MR7WLOqzAXd84j7TSIw3J+f2WutonawTW42oabR8jr5X8rUaXgsHy9ygdIT9wLuBalM0Q
8MDw/pMyh+PjSg7MEk0c5XU7M3/h+F+XpbILqNmiSZpOsLm1h2pvLPTJwFdNd25uhTRK0mzj+Q+L
/dZihpWm1JON5svp2pBpp6CUxevIP5OdraPJg+fjTAIbpMsrb7yiZwJfqcAYrAffWwC6CTOtBHxe
qgkSvX4Sm3Mdi5+brRyDUYl2inoqqzszOgaIhY8bxdPgicM5x9+y2+iDkd+gmPN4K6XUuMuRNFbx
S3THv0TNUipXrL/CMhbFzpM57O0MyMIcklGbqAapj86OR4yPOg8zpBH/7tCxg7lJCMmL+vh6KFJ0
djQFTQSzVNiUW8SrdbVSY4Jq0xxHkSU00H99ynN58tCga6eDdWm295M3ytblfF0smDpoBDy8ekcl
K79Dy4kLAg72zitbETrHZd4GS15D/ARAZmGRVVys/w55RKBt0Extd1gAoYbvgK2KjHXTMEELUI7l
/XfFikpVLxwUI1ybXH+qXKLsIcnk0hlFUNkuOP34NneqCZoIxW8AuygYX2F813VL+KLnbHJb/TK0
zdXKNAxC3akUVtJ/lcemtEuEuCwA8VrORLexKCazxhlZCagYZoCXObH5KcXEKMqfcIUTgLDRhTa6
BIS7Qq/VP+UF7BU8mIYhtHwUUFaJSuAYSZu13ald37uNqXH8hS6g8qdd2mVQnxSALlfkSC8ugX3X
NrNawPH3hdVJ50cVX8wnfCnad3UEkqBSnFyVXzkIEdBmS3exHOk+ASizpSQTbxZ8qADfhM/hdZTB
nM18mGMM8jzL5Jv1gUkjoBFxOHlFVTCbwkDJTwCxHd6Yif2Xe3SA1snGKEGYIbABRT5tnRVBHOrp
ZcNTfdWrcpAObmcTnNlyLlQ+FSI7/nMR3OjEIG27k+KVGchIoTFecNpdrMhlGV7dMMZT0fGTJOh7
IGFSd5/J6wyNFLtXvSXybXxyd6JXIdRVrH8Ye3IEs3iha/agbY5n0CUronLnwGptzj+onRvjGSV0
1QxunRpBgYeGggCYcJTKKohAU0gVgEj3DpA3EU0bn1L0/P0GorNcwSHx1v/tDowaGxVFhcg1Z7RW
p0/63e697kv7FzvqdziTQaTEpaUFLekZvVziD7TvI7LY310foPUPq2+rAEkoq4QP7CC7tTCb8RLq
fH+Q/qtSr7EqSj3ebW/YpS9x0b9qveLC3LHUWX5HpaNaXeqAcCcsWhZQbVAEBOHLWlFogBhCo5RB
BqPmv/Z6pARl5nrXnTgsnqjdq6fSY4ktF8/rZcOMCUM5T+cXxGk6wXxu2JY/hCjpqEEUcgDcyY6q
Psc99FCgCZUETGDSdDefPR+tmXdVYV13FuF96QctS64QgPKLbseUHvG1ANFQQ7g4sEYamjaiBZGJ
mRW6rT7qaBFYMWSRajOvHRUNOUWh6j4nWwmisuxyE1jTTLbdaiNEOC1nqL/TxSnvEOJ8BrRdEdkD
e227DOYR5CBf3UOSDxRSW3P1owABPi6SbDnwNS30vqAxrARwahjIbXMvMxtqVaoqfIR5K0ylRxo7
oSiRkJQujNzfeLbVIavgggqM6I1I2iFWKlaV2ZFujkaCWdmyzYVq18oiNGhcnaeqbWhJ19/eVlF3
/TpOZPJ3NSPXW5M4GgKIc1sE8UqYUPD5OXZxC2R+WfqNwCRv49ZBsRwZshNg/zNZINifL60PkMo4
lAiVlbAeKQar4ERi+Z4NgDU7x3xtvsJcpNLuImsYvnwao8+x6N9bzxz0rfAUeMObJTwxNYUSXcnO
3X+mDzJ3Vtcs1rykvpVYnKrmbZ8iI2tzafRrROeCgJJUI6aEMIDHpj5r148iSKYtUM4jMUfbT2+V
PyUUjzzjK9TfxpCSp+SAztKmwj4P35ivqwfjW01nnLm2DYqVzxOuhI6toh8Jmep2e6y29Fp5gwIb
HiSjfQ5RIwG7GeDj7JgUuk6RRIz+JajJdTaR2Bjg+f0H1wRLnpsTMfvHJHJVfRTnW4AHUqajtV4W
DEcBtUvpDCj1XCPYspZPVNRtO57LGRntfi3aN+WYHEow4ODo05pucllKFw6pUao4/r6MlV8vhuf3
NjfP1ReOXel+UMDWYqum2B3zv06oZejV2h+FXtNpGcQi13ZXRC76c4jJ8kO5VKZGppTp1TPjz2ct
+KLUUVhoLiz4AJK572kiQxmqFJXjjycpy9UC5cKJiiHCtbWxyk8Civa5Rt5pzhIDixcHgyfmtWPl
4V6IEd0z0R7OkUtdlApg9H1zKJO9XXll5kzCFeMWS5rKmQu3MnGr4lLNpzRzdMI+O6jqysRB/f/O
YwaJUdEGJljeF3IsbbyiLhUwphBTZD2P6gc6VgbzkuTHHTU1ZjW+mX5AvTZ2xlgJlxnxc12JHPRe
mQ9FHWDJ0GvmZ0XGE4CzuFnXZtPy/F2xgxQftipkptMzi2Nq1BDJ7tKFcZ81bWVLMxgwh9raes6U
ifL/XRggmRk0ejxFpdXsJTIbqQQw3uZOdGYdwdX3u1lnv7zIi85U6MiOg0cJJ+m5k9lelm25Kr2l
CBo6gDEVDCT4ehS621QuoYfc4V+L3ic3aCkKh4bQ6oM5NzCHpsojhhSa2GMpD9CQmh+saW9XoSut
zLa9JmEtQgN6ROK9Sm+Hykeme+ZItsjAtLzHKgLFiyDJywtulhvH2jgLpuQCBCG9I2v6ALDYNw2F
t4LeRbeqMUHC3Nqq3VzoP54nooG35Zh86pAHv2MyGZPb52hFDC98H/eB7AB1hnW6GRGOMrQNS8xY
fOhc+5RTCtrMQAyefDzPwO2XsFR/e+CiCmQwjyCqoT86eQ7sD3HL5//q7wmDWCkzE9Vd8VFhEqU4
/BFylQfY2tSprtoiWjnZG7KA2BBDVpgA4LMyfoqMPZDQmv6cZDKce0z/598DeGo1HJaYZ1j6ngTV
KXDCwzs+W9T3/7SFuKOYbG7/cfFv0DGlaNYx10qyZVa4FHt/T11kKVbTFVaYIBwzJIZCJRChTECX
MQd29yuu+9LAKbpj4qGCkQjgiGBrJBVzyhhnssNMkfD6eP2TeSxibTjYf6A6hWzqDhZ6Vwb01Tau
yeejScqMbB59jAI+9pBYvHCuDmaw8iGKRhwMXvXOtM4IL96BKcZWzMI2qXMvf95UDjyFH6BOPy9W
sAtjIVv/eGYBFYo1AVEDVIvz/BEb7yr5U4+j5Wm4RBhXGuNe3lAh7ntQMNdA9AK44siNrT+jHCTa
vrW0xAVOA9GXMh8RJGqGrwkBeLf5UnSXP6ZqThC47SrzMDHNVGFbZNSLnIet0q3592nXXNFhOejB
TK2VD4p7W5w1vTuxaHZYXCQbOGR/lMW8yOAlzzAmqdb3EBCvFOj16o7+LYwSihSEgaEZsg+RcBnJ
vRDqU3UHdr5/PQgn1omucR52AtIJi8lurjQjdSwZiPjfLuTjXdarrhtQTtszgDiCW2Mil29skPvm
ectDkGMhy3CcOGHnFFUBm78Mi8/jFGFp0aPUt8hEI1WPySWvHiZLDcKNliVsXOnh59HRhRe3kNT8
qWHID8weDOG9pLZnMpvlr6HITsaK3fRebmzRZP1O31S4wgyNO0RQj3Y+eIpE0VdPp9ht9Oi8ICTw
5CRaJc+jq+YIkX7fNF5LHvNN98R5oB8ROfkUIZ7QMlDL9FRYymgd9tJQToQhvSU7lddd2PtBUMwY
iRKOKSAqwsOjsvOZR3iY6H0JVXNK1bHCRhhr38L/9GLkAo7pCVG9nnkO4u7oQYl1pEWY0Lrjvll3
CdcbHDlNXfxYvAgT9wdSCtpf7g8usEMe6o827AGv4tTdRwI3Gg1WFAqUwa4W2WShwGZikM8KhUL7
gDpz41aG7r6D2P1WK3D4UHOchIoBEJxLkBmN1TQD2xQCa0pFyn5gAN8EvNIDWecapIRXdhshWc+2
/x/lhoYKv0r/OnCX736gtkyERElj9TMNE7cQODA20v7Aunu8cGYf+iarvwJ2MqHbvpaOR6eiS5IZ
9wTYUaKQmfEarvZjfwbQGSXF38FAsO3eV7TSHTqEUeGCUvoMBiQ1TJbktn0Vggpq9PITsTB5e/QZ
9j8SZ8t2mpZ6F1aGXRN3QmEUH89kqkc6bEnHyAMaV8QrSOjnDX4uJqStlJm8Ry8a4uKRK3rQSUE4
5GyC8nUD49YyiQ/pkboWVR6PDUto4Yo/6InXhS3Zl391AY/lUUNrgOVojQYZascgOXJfAq/1smbK
WRXSG3EdLNbMx7YTTg9VRCfBAmcUPkFRtIt3jZd9ukWOIfSRBtHridaIhfJUkmDiBCMGd4lmNfm6
ZZ35RtyJGaFTAp+vOf/rs51DGvnBe6cT96C9VlXShO+SXZoanLKIXbtaZqzyEjHwPmgjq2kIsgKK
etE2tfN0kCN3XfTAZ7YPfc5E7/h2O5E00PK0lbRQkuDz2pK2vuyutH5SM9yCEQStjwWOxuA0OVwp
BoZ9zKmUCax/L/pXp9J0YdwBLHFTEyioWriB2kru8TZx3QFqYbgCrNd7s4evRc/8ddh0e1phF9um
9yNpQ7vSR/4l8uoYtMphEvXRGabXGfxt5AD7bEkLxI3jnLq2CMhGNcdzF/DYeEqpHleDYf+Y08MX
co4SttFDaHMuA0jfSaY5hwQdLCxJdxUTH/hmlxdaPFxac0ih+IwADKNTgL187sCtaBuRB+rFSGQj
yFp4sakuwz3V86PPolVU7BWC2wl3tvTgABoyT9Hg1ecrl2Qctiu1OP198gHzQHbJbNC5X85Dszi5
HhevvpKIUcCyy9hd3y+Xy+DZ63TyITTNyfq0v9bYJOyDIFpVddjp96wL6PtBayX5kBPiuh5wQyOM
VeBMKAop3d++4V4dcdhUUcK+LyCrfr0oEc5njuOP65wvNi4VntXdwmF9hLihdxYt9zCmvaNbLuJa
LZacnGe+Bq/ifViZ+AKV/9Th7HFeMCERaJcv/uM0t1DGrCU9OSDJPJ5WQebLcPIpywOkTXZVFZ97
uFOs8iG4FzWTJL4CjrY1ZothUtPCT+rdiX+mm2Eyj/rUqyruygt3HcbjcsaTjGdNkMJF07Bm4Aln
sWgJPAI06SspVm+yaLCA0quFN9f1QBOyMAZhN3i0wB4sWV+RaS3AwxBTOtUMfYLRZkLVmMl0s/WV
M/1ZqOFgRyG7wNv0nN6Jvr1jPZ6QTgJ4bJP3nNyvsUaaCl4bRKORWMrLyAde/M5GD5z1sZ3SKGr9
i2xbKgogNSeyi36LwFV5iR4ntPxRLvYEhqugt0WNiIW829vONZr4Eh9DqAVrNzipxFpgJmt89sMM
R4uot7XFwqfD9FLgigKQw9w+x89XzKgMj6HydntzFnhJU+DvsNwfFoKp0MqyM7JvDdb7UREjy/ZF
Cr2Pi8U40uleTJUsC8TX66YpEGS5pp0zpmLr3gK4haZauWN7iqMyeOtQEeMjMldcykhwSZI/JP5x
tkdzZIsA3VEnH8GdRPRpoFy4FXy/6cfCegt+Y24wsmGBbHKmYBSjaL26Fvxs2R0erWyvNjdif1Wy
2ALpetsXLwGoo+pqWgeUGEwASufBlBeMqlERXXipBZfJUBrjpKHX01EZyBEFy7/uufk2znlFJFWL
Sb9eLarTfsqk4grUlizmYedf4M+iElRYyz2RlsJlgdJNj4G2+Se9aWbNsNAdI0ctmmDQrKweewvZ
R3ngUpBJinJIqZxtVBSpWwmu4+OLHTHjvpJ8HyNIerXrEZ6ZHwvPPHq8RtTHkDZP7Ea2cLiQSVxL
8dYraXSoR8dQqINrPnjntfWS5yzwB1Xwn4he3N4G36ZI0CIkj8jKGFku+QfE9GLMZc01hQyVVPiV
yi8m0NLaDgNzsq6aGkPbs1niLTsrNIQKe+ZXygcvCKQvkGUQD6t0Be1mJKyZLI0+cGO7ZarO29qz
eBFqLcQK9F+aNnOgqnqWsAFzZSjo/hqD6k3c94spYsQDAXdHWka6AQUruQRHvEwWF+R7hdJrKQf5
nRQuNViF8XTRWsms3rkjq26z0AsAGp73NcNA5htARF7glRsW6FJXlP3ZhMCsOjkKMx3drcvJMBpC
1NATf9Sq5mwOipGUlZv674+OgXb1Otc3crr10+wIIkEE6r/xk3vIOdWayb9jeU8jtyhrXRsZfdTd
Onau34xWqVNjPFH9I6sPd5NCP4v4S+pzd6C/mkrYGUobmajKK0bq1KnqHegZk6p8ZVCvL9ncuL7E
XC/VeratdFg1eO7lvjUA+ZJrIWOqYXMA9GkKtVbFkaOiGhYCXZ9RFqBz+WTDUPnKFY8MjVWHA5mN
eQUF2r5jOfdSbCoQ6+/0BnINuqng+mIrx6ucheqf+Jd1kac6WToqRfZNqXXdzGvg92WzYEOGlHA0
psaMyv5XD75wyumtHvmIxHHNHAT18hYTNsmuOR21xhy+kZNsTY6jWT4WgRk2ZzIZMbSofaaNP0A3
8RfBBBWwf8EkRA5IYk9fPKZEKeua0rgthc2NgT8lq5Du23ZJ8CCn6OhZZRgYT1/hwIuBAW6wZan8
tMSoGqjRcoq70ySRiWzrIv7MtfS8vm2A//KjtMIDoqYfnprrWBFy6SlkqIa1hwG1h1FRaZCbPUZA
AK6UUGdhaE7QTWsMIX77QNLuc098AvLnHN5iMe/gYYbxGweCFM3FzDewnpxjk82iGDKOyxe4paKN
k/iIfEGVE7NcR4UI+zykGFKvOIBl646TIxuEo03UIH0UrAiaAOHDLp3yC9a4EjvjWiQp3+Wps23y
efHoQ6CP7OsoXtQvsQeCdoc/91Dz6wMaTb1lzsXbw8Pdnc1xUbt4dqxYOCULbvCmz6gTP8CYeySK
XDqIyBnAHbpr9gRKucCpHS1bl7ss0agASWJLbEobfRLkVTT6S7xs0MkrUrD3+VsYJypcw9hFd2vy
tzCx3rIBX4aCX8OKACkHTuNisbNvo57uxyu3JmSUYx1y5Sdo4uoRNAUuJhC0rJa/1n6SG2FmsVcx
dTKqf7PAtK3IYoNQ3ZdMeHq4GFvzkFiWoLlGG7Wo8T1jhGKqoTMBZmRop1/0wPC3aoHERRHZUrDx
BcC7tyVTc+jy3+BMPyuyMkMe96BzSM2Zwyb3j8xWoBZaW3Ra7H4VjF6QuD0NOTjn11O/u6Cs4S8Z
XJiFGW/gmC3B/C+Vky3rtSBMXv/py4A3tnO6fPg0b/G1VDXHB+8QteMax53FNcK09S4Gca0QtAtJ
ltQ/YvjyhdzqAurlmjgRPOlB8Be0wmBZYXUHkplnKOqHbKfxauBAuaJUyE45mGPISUXT4vpnBR6K
Nf6mOGSHGDG7MLPeK/kzfDEtXA+KlgPzpJ0sy5J9WB/cBvI+hAQXyBnrTwllKSnB48xV3J9wFgb8
fvdhjuAhelXyZk0L1uFTsYlkIrA4WmuP4dMTsUoUREAQJKxXbbmiX3h4g8HkFSdB9R48CMQuodkW
MExML6R30ds7mCejX5AuOJOx8DLaHR6NP4CdAy+OZc8dczy9rGn/0Zh3J+Yq0FW07Y8M1ArilEsS
v2TvSNAcuFPGeO7SPUrRRPynFnqEq3XYxLLZITW6u6za6IUxF+uOE2hhMJqnqGfUqiOjLj5OoSK0
64poPpNgXHPm9N81ntp3eY+Eb63XblidmeeK0rv1Z0SaMZXXFHAchgXeF/STngrmW0tOd6IYIhJA
wveSFSEThPQezoMmWkC/urOKnH/x/SG6BWxUq+fWkpMP7/XLI+f1TIVkwU29lYA3YB0bwGvjELis
l4TRUFQUA93Qt8RWUA1PzoZdzwms2R3fmBz5CkYNQpyoclNHDBkSdsXTNEnqYKVviaNjvwrL6DR2
LOPR2IZg/xwtk85SwuVlPWgwgGiFC43mL2y19fA92KVA8X7ropZ65hzKxwJjEUl00SofuDFTP+9/
sf6ZGlt96irqWCEyZrjlgxMSSISw9YduRlHk8LFmfmIxoP7peuwfad1kNbBfONl4br+2j9CXJAzX
iSxu+X3eobLLZCheihwrop728hLMGcRINqMoYRHFz9hn6lxClHPcCuPeUFNRYpLfIIvWNbYcw76I
3MgbkijgT5Uq8tIEAZtm/qI/3rr8mkCfRWbNVcBsS55V8UMLZ9GyNeH910jhLpOwkuEftj9Z937O
9hpjX7Bj/tNnZoH1p8unoVGGmBO0xTix5lgbov4cmqO0GQ+8LHT92yf78st6JVPp5dQa7AHL6exl
LHCsP4aB5gGrbUCzbNObiKG8hzOUQ+jzjeaJkzWWQvMcdXsKAF+EKndFLmYWQ6xHj7nSJmXjz6gk
oW/FW6r8BHZL9/2rAfriZ5lV5zlZwER8bH0r3KORDGrySJoReoPQWStzaXIK+4gMlmSmS7+NiKSj
7Y850eAUxVszOxU4jhP1vNO5Qj9P2NZRGnxzkH0wox40yeIyX0VZjmMvAA36olZmCww0/QXL6Zyh
jPvPvKgNBciqPDJFiYWFBXcvTiVDIAvkSxaCstOLvGEpweCzErNsXLz9rnJeI3nOFQZZdLhrt0BK
dvnfX7YCgHBYcNdl2cVeFVjJhabfVp2co4//GLb+Al8xXtdCZsmPRZLWpb2jv3ElSEIfgumfjbaH
SVWZaQTHngpxW7w4b5NJe+pUSNDWhq45cQcqd15LCngTcFEmoY1AMfxh37EzMeYved8ptGWtar7C
zykqYvmWh12enwyVmmaP+dRTOykd77JoZfIZcqtK1zLuAiQEf2M7/UECRJzbhJKj+fxTgAbmbvhb
Ljc+3zMNu58D5nLuCfUmtLUTmlGIIC3ggcow4dERV1DnkFDu1aj+u3B57YEgcXQ8umnEZ69ScFBf
7PsulTpaB9heLSuFu+fhzMTz3AvB/A4kL7mV2gR9f4ey+qTMvNIBLvwN30C4XVdy/Zc6IzAp0whQ
7DmotEDNG8v64sW+tKbouKA/hx62+/qy6PLKT8SVtKP8KpITwkcKcqmvYnrjUNpkwcRZKPDrCyMQ
Tv1bi49tPlCMF0DK0f0Elc1f/XdDXwFlR1rWTZZnjqITV8dVnEDSn8rqj3b/uksG7CD9m7BI/Y5S
Wq9x8mVK0tTwjI1ml0bW38jr5bE0Eb/EVJJLOO3riLR9J9Yhp16eBv8wrHR/nxXy9k+BniSiQmqg
taAQuqgJ9n0N4fKtp46S9dOvbVYHC/YlIKhnlI3j7GT1WTYDHSrIA4ZESt7AcD2mSfFSxjkaabDe
WBEnjOj2WxsOWDgVVvIepMyqFhnz3n1m3Eu+Yh3uFdRdfwQC4eDQk+sPvvAl2F9YA0hEiMjg1b46
NU1AGuXZoURV+JSwsLb0a4CQ992fHuVABb5oquOqq5uHnJhpMBL+obHokh9rN5ZO17qPhcsgtId+
uE2lZ14lwfnMezD2HAadtM2NfmudGLlj5uWiZhVh5uxEBTu8DSwW8VRctIS1BhPDblSsPSF3UjJ6
D83K7A7Qyx15b+85cWSBxwZHqQKTKSSANYdhYC+fFUZdfdDHLkGfLwxLtge9BoF4vhc5M1nxYlPr
htB06pDljovXIr7KDIhfFwcRltoLOc0noQigSYRYYkZj0TWwi1CAgd1nxNMZJwOu0hd4CvYeLn6R
V/2FQdxQaT51y/2d8r8PGub/1l+Nl09cw9udsRY2jQVdLK93xdwQj9NixTFYMSGx8rG5svwwdkeb
Y/yKLW7LBJIHTjAvJfr/XKT7NX3dRbKhXbL0DDBH4yMGrflDqRaPdVa9mKy6maeN0WBKkfUNQwO6
eGER/rKZRCfyArPIYhX0Xe+bsEi3+jbfypsxpeWbvdgzjS/qaG2sA4oei90Sp1BVz5U/bdQia5xS
ujzxPB8t5f0TjkSRmcdtsVQ/Lpg6o+Ma0j2aWLnBCBUnhD5TFB3lPjGnT3pfODvpHCBxjmApxiv2
f1O31Rd0yfB495HQvqxgb578kfH9ixd8NnmDhIZxvytEVo6Mt5feiYdIti1LY99G1FUGZy4BJPm/
J4nWpbNuo/brVflJFf7v8sM0/hLLIRQOMRqouGCJVGGCVzGW7Buyh49A4XCVGjt5t4kOoBxzhf9b
dNr83d0kD8qjxyChmugjooyWhHeV084lK6RMR6hbFl21UVj3Qe6GYDb7oedsboion/CHRMwBJUZG
LHEtKQf0c/LMpdhRKCii7Au4xqF8xvLspaUkXBUvNQD37thD2PFzVCt2dMNuku2B6ezmkZ1qYC4o
HB4yLhrC/z8ARoTi1DJSeYUutU1PLji8MiKgIS4fKgVKpjJWILcRvrdCm5gSK+i00xov4bv4AqJW
4SHMz/WpfCV2sEswkRzuXCsK37jtXWzJXdFI1K9v8ELC2HWmpN3M7IhVFe3zecI7YngiqZYJ/TvG
k8rAbN8e8CLV3jf0gIY+SSNhe3dmAyrJD8vw4BBiL4x7Y7s+5LPHJssBCAYiLF/SPuTx9XKxZBBU
xDsE/6EJFs6ziZlR4cTQ2e6q8V6f2FnWpJlCu3DHGePLNjve3kr937IkET1FID0Rts/bByFVibMO
YNFmWdiWdxxHpEI6VPFAUJSt7FMPZSMcvoqPgIRWJbrW4pvJ0Z0TrjmORgCYWm/LjKwrZDaIYBFA
yqiZWQa1q6FJw6KBH7OyZY0B55PtBXCgOqba7/02Nv6/hqpU9dr1bNQIsGEwi5lMfTDBfTrJP6up
Wb4G4XX1km3sKnyECCus8rMCtIj0bRTZkpAz9TVn4fulF1xEVLSkONADKsRSKOc27tR0gmUYKuCg
YbkkLkA+oxLeC+jI8YFJDrvMKpkTK9izDKev+UTYqD5KNTwppv1KDVG0o0tvzVmmXB781VZ79OVZ
lDe1+l/O0lNsuiB8TAiEMBG2HtgO7TeBHgxH1zT+MZ5ClL6BNvCLNnbyV8d019NWrDZH8zMZ8KUI
QpXTiaKVDZMSlCQ0CFYESbF7OO3BHvLdwP4szlOmYkATS3C6YJa6wNM29OSw/n5NdbXZYTiPpjND
gNA3DwLdOHspyCUl6NidGthTrT0Wg6sEWAUDxOxu9S46cNdzRIBjCQDN7iZH8oK5bzmvL68Vc0RF
9GNAPVT2mBaFWz0PY6DZdtYBjSeFv6M1E5zooQQKNnJCDoYJv8zbO+YSco+EkA6AD9fmecSWpupJ
NtzPn4w7G/83Wr4j+CljZ4m+3aR+HRDk5HrahnPOwEqUamYu+3oM2D6Usrm2yVwMWsVJV6w1k3Qr
GutkxF2zx+z8r1aZaRLpd/JEkTte+6XX+Khm/WoTK5Ow31+mbry7fxcmUzxtNMXgw7WrTAHTYj25
M1OcF7ib07d3QTP+w0dhb7yrDM53Gx1Y5+ExIsVrW0gfcCFKBzOs3fYxcmijSp03KkrY0xD0Qgxg
ar8BCj9fkz0vPaCFj4T1Bf3Qx7RW/2fGx17guHxB7zHD0Qw9dvh8YAivMU/hWXJgBFrbx5Kn6ZGw
6ALhqCYWnnh425yDGctkADUg5xzUlKka9MEcsJt1vdnWKfG1XUoHXoEBNORRJBUGM2uSxVOP29Ma
bER82mFeL5qQfI12ECdxckIaQqGk37zOUN1ArUO1BJzY8go1154JuUV8Xk1Wp4qW9yaogvuxUyFT
ei/rlfQ11N/czT4ZAU86hQV/z8KMQjPVxGmpKhwk4cq/gzH2doPJ+n3oKVuAmKwFTbNB1Q4nsIRb
5o0uYoxVDI6H9QoQQ4UOZQpvsTNcj2RjxgOj0oHcwxqdqfI84gVlZGjDbgMTUFp4nUecLGxZmNJY
MezO8hxWDqvdQWFsUiMmtdRRx8t930RjGr/jfpeXXQwmfgZfk9LBaHUHfONeVt8VXJoMHKnbO6eb
MQ79qXW9aP8IiJ6/83la44eHG+hJaE/mMV2m1XhKO37cmm3lDvfTLUp8VYRn/g2C20BaFhaWADUR
JEAE9KtnhvzIV9M1YnMZJ3iLqtN0Xv9kUfGsGQpQ9VBBM+6Zilnpd3tbed7dC7jY8PLQGReMu1Hz
ak66yLg1yZLR1S9Bg45iYl5XA2L+NRb7qZJ9UTZwX24TQU+0y0PwBTQQxscdnIhkfYC+GuJgMmRb
dbS6lGBKzoK6WSPlTafUsp/Vtb26RvwP1ZMAAY3NB0FNKvuBUMxeqL+e+zhL2PUQ9A7/V+qav4/k
wXn5jyw++04T/Bvc82ZrdsS/zFYkQfE7O/sgVPVltfdS6u5TKUxeO4m2J04qN1oVeF+zNGkCx0d2
l113cOXb9Qz7X7NOnjfrrkAAj5CjK+QCu8sJJncHqagids0uC0/l5OdDXzHvfmsIVdbqcLclH/1e
drVyPyVj9y+XIi7dqkP5H03rL7BS7AP6WxzIOEDc8rw22YB6B/rxqsufYYPIuZNc3DAdFR6S1aJ2
1TpiDRpU+bWCAfqgwSOLAc7MZR1IF4Ahj0+tpwsXEoLILgRkyDBcAHCKW9HDUVyFes+7YOwdnDYg
m847/yVn2OvtB4qvkBqL3nKkPts9QNudmA1vegS5O3aeGSUGiuxRrD+7Aa0jOUN7FPyTQZXn1YGq
Fk0j9YZyqG88WauaUmqdfrWYq5WyWRSsuJ3oLaz15EwoDJZC7+tgh2AvVOKWhw/VS6OvKo0tIyL2
pilg8/Ef3k8eEceHux0znmG++/bUVSJYaf+lGiD80/Egs6+SunuioKCcYF9WZoee44ak3O7tSNYI
VS6+gTlcBUjwQdHbUt7MVM1bhQQkgUQmNwTRV72a7x7oBOv4w02BuccYMQ7aET70zx0JF7BaITDA
Fri9CchQUNYO7TlzZAezBw1r4OuoNFRrODDWJ1l75HYRMqry2/Aqneo078rtiGdrWV3aHjSrmUzu
YS+v2/MedljKZsq/AN2cTCs6wqKfsXmRkqihaCNMFeTm5IS3AvzJSRo4KClrujRJpHIV1C2P9zGy
L52xguKSgAKX7Kdh2wMAuLIpqgnFH/zD6LjqL9Qlaf9vo0UqWHCSIFfER6BBJbra+ZdOPBWZNUcT
2vnqKp6HYgPQOtI7f2bmsDnbAo9pm6bbft8+TQxq/lPM5EdazjnUVHHf6vAszkF/H6lPovyRbgeA
68ukYS9pQqA24/lvG6I21WczxCPT8yrwYtMpaAFcPSZSAnQeFTnkUC8x8sMVEqkyn9KjsTXJNo7g
zYlYkn1sb+shBjTkcormO7wgC3haTCKxVYJKCsZNgj9SNRAYBa8wTRkmA5CGSp4GLJRbZgqnfygQ
PHVpyKNUNXOeOXEGk3RgmJASrvFTHnfc0d/r/ubIl7VAIGJVT5+OfThMWtesPGKZsGtoe53IIj+x
8rGOSi/YdoVQ3DUywYyJQZ8XFhvt04T0Ve0cCOwHpblJrUHt/UfSbdFEzlryEtT2Tra7Np02nknG
sBFJbY2dESBNh4XNYlQHnybUdRlYbSeeL4g+5fgs8FXcEhGVXU0hfvXdO2tP3sNAF8Zl++Xblppl
Ebndcq9dr65C1Cbnl02UBY7iI3JqKjJ9Jjju48jYU2KgEljZA88BNWyy11KLnNifPiZDa0I8tYTk
PTr0ixx6HZW73khraXH011IpJwAqDPI39L6eF3LzHPhfT8aElOqcdtI7VhPaOkiFvNsJiY0vFdHx
OOAWWzHcBieDPMwb5RNtKXViZs5fZRPqvahimagGj+w3mDA9hBVlY3dmywy2lAylV7KPxndPcxQ0
lZH6At8whbysyQnump0rIBKngQQVotAECmyMcWYaDtvXjdTe0vwZJ4XXToAuivEBzvnfZlH7HXf9
9vklkLe7kaLkv0kZkdjrdKBsBla4RaoBeBxLQGpEoNhXCZ3atRaXqBDOE5gQjVCv+x2dDxANrHqo
aq43an5fIXJ2/HdF8xOehqCh1JqszTaBeG6qvMs9d8p8GsSjKlD0bgEj2/6YAtHUf9EX5CR8WGQ8
MZzmLLfwUggcHWXUH3qFm3ahwf2u+tSdNYV//Kw73y3dfYbvB5PW4/3ab23swZYtsS/bTgqaB5LU
qHL208QjPlUMjsUeZbC5Qg/eGlO0k9L5gUB8VFIoHCLIsd+94Q7h+mOSUCLzCHXS1gxDOm/RNx+j
z69NtwrtoT8jZHG9lBGwDh+G2Yb8qkznAlz77nLKjpNJDRRufxVBpYUS7R73I3OmBlxbLNCmLTIw
zillxn2sIPggoJwP71V734XCSfFrY/siYFpfwqwpwP3Y0/r9wg2wcKPHaDEulBde1FmVb162aJjB
/3bCgCCQKu+C7bRj6zDtNJdakIRJJizAf+QHG4AIpxtrgZ68C3uLK31OcfvpdOpLnA2wYKBeUZXA
1Bm6fkhDyY6GdDZDSielpsZ7kpcHEpwHmwCuDZfRepoNpRIXsg18OEmmisGfSyS1NCT+HDn7CZ//
TK3aXqyaXVk4CoZoyXFwQQkuY9zU8ZUTDNpS0mTVauRB1m4Ev1UZ6q5QA68NAFwdOwx76O2RogOG
mVAokOh94P0E0vROfJ64Pyuv5KRJSJteSqF06dZKV7wOTVcBpUKMtvPAbPyhSul2C4BX/QkRieIJ
9I+WnbQ37lpe75RhQQI1Sy/uEhGJwudYJ5nievyPR+iKSzS2BhGiSmUQUGd/9ssXN6s/gIjJzVaG
AquYAfwokpdqvRS+CYZ38GqOL2sYxqnGFmUPgyRAPUoyaBH9ZmnS/uZ5vTAontQEq6y7x6AwoxzK
uaXPXrMvUbxjpi8SBeJbAUOIiqpB37NnFkIQjCRDodSZm3aYdtM6ucitCcYtqYnCvLIGrB2kmHN6
h+0oIt2i+AqnUIfTQUSBCj4lFUZl9MHDu3nDSgMG+f3aQ+pSAvDCZ6FKgt4BpLmW31InXIXdFun+
GboJ+ebgf8KYWbHJ3v9vL0cU16pOCtKtnLRsaK+hLf4pHIApJ5cPKnbwWVsMmfrtIoX/WU20Ybiz
Tf2HAz5eGGilYyXdL35G48rpgFLkaw6nbeyxFFSHcYTvhk44c5ZsWLNyY2mW4swUTTCRr80Vssra
jSZU7egar8w00gZM+xB5rEKuraRQ78eZ1kF1+hWIAC3fbat0Y80Ulj6BnqcyElqyby6Ywr3qgk2Y
vfT8J9GDZ6ctMqGVfFl6ZgT6DY0f/umYlXi3yrNcvT9lRAimI100yyI4D63yj2cDSdB6eUmoVFHa
togJWHhT1Yfs4dlpOuiyAs80XMpwrvsigWm8wiVX6WCFFZyzh45BM1osAPsr+/bdBRpGnJ7zftpx
3eCbRR7zu17/4BidbcSzn7vf44qehMyWRGKhiULvD/GgkR0m4aLf63R3hXFgzYROuVxGaiZRkOvX
sZfV5/Y7ZsG5DjgiPwzFJDBn+IB9y5UV5XBiALxroPzNgSnK+ne4vpjIxcLMlbpdPsLV63bdIjM6
qUS1SI3boIepHFPt5ujYbhmIRd9FYk/GgV8Hj777jMpjPKWH5Ds/Jx95o3/gxMIqypngr/LAPcoj
LqnJSgtADAQN5ByMQoj+PDZe14bmevQQMtzRAYbWC7Lhva69z6lFYrAvRKZshgkTvcmswgysTC3j
8ReOiLaBPNYtmV69lgWS5Fh2v05nDoHKThxndMTLXJ94ZgdFoFuCP0dIzkH3Vhp/Z68gNO60Z9pH
hiNv4pcE9VZCQ7EbBK62TB0BaNObdw0kNFsf7oVk0p4pNbWg7P67hyMJSgQEkLI5WgMuXJYKF1rB
qCQzsYa34rVHxWqerw11EeWfpUIL856WS6HiBWOyaUYukszGTByxYaUefcx9ZsCpCZSgAp/N6/3t
fkA9ia2RFjkVOf/QH8+plYKvibGWdEtiGkVIuCgFs2jsMYP2/xiNkmB++Pm+LyWA66MPk/2xi/ji
m5Ke279vnr5D6u/q9ZhmMoh8Rd7lOCeEr2yR2KIBR0TFIBeZXeM7WeKUmPOrdUEVx3rbJxrNiUp8
Pv7kM/YDbT42Nb6rcYy0rY/rHXa2PmTUdCVJPuRkNYTaA9yYRB7brD6XudPuLK66MLXldhBxwJIY
POIGki2KoNmnu5j8niINoKVlDMYLNYIspIR+PqAe7SL6ZGkgVUdBjDeKtPRlWh9Pq3p/uup6H3co
CqcpYudFyneklJBeXsxugzErX0lMcXZbi1tZfhv+mWwlSIZAEy3EV1eOPWwolQgEn6yShpiEdKSX
cVcRGHS7bdCOJGxwtKeWLqUuEw+7Y/Gjc2RyMPxIWHeKvvFhyASrldjgsAEsTebej/IimYJduYnp
EXq1s6ZNkprH5ZJN3P46sJIqEf69PqsM80ttPn855Nota+IBfFnEB0r9PLnCd65e4os1AGxrF5tg
f7r6WOAAHFrSjmKu8fwYqG0yFB9/nN6p+ItR6AckKi8v+gfl0DhQU2yTOlNxXVXcT35c3IL/1k99
mrnTkEQ2BcMXSnZ+HULFlL54G0ShJoPewG6ZhtkS/0oS2ErUd670kI+14ERS4ANx9YrajoRled0Z
bmSfQeKyMP6STmwyRmCSZFONCQRVwwZrKAUDUIYn9i1FiVZYJ7rP6fIxB+3Wf0HsnQWh0NBnJcxZ
sSzHFnEl+4gI3da44Lksa8zFysRI+Vc/o8EAFkns0j8LwTorHOh0ASVduwesU8DBCjZZD0sZgpXP
c/xyKUC+zR8bzJ96zG4+QX9RAxoeRfDMEpROZ8OGGOmqeWtUfDc27VqYr/q5SDMS7rHpijc1rJN9
zLPjhislTsyL5myMJi+j/I2arLEoQVmKWnEbXSKp4PdmIWRSDfn8uNo4bkSefS2//wlSOWLUTUzi
idyz/wAwiecu368gqCjBsNQOdAtr62HZDPhzjm9KT/YjOehvxpj2gThe3g2cGlVWFpIAHDlvub6/
fKesfMInvIpOZmWG8xXpGRh/HqyFENZIda5b+9B4e/Hc96r4fPRQWxyR7dJKiV6cZ75vAfBnm0ju
xwqFMug8FO0p1R52lWFYG7l9M1jpNIUNkJ6kXu1JIrHFblbrowe++WL8x2xHStQ2fd7CVvmGg8lf
bjkADP0Bfa4TvLCrfcFQG2c5KfwpEsSSEI/P1gj/bdL+p7Flo02qCpluMuoAiT7f04KvyXBpV8Co
I0YaJUCUWGywsqYpWYmBECmpESoNXS/Y4YNzCHHqV8j40u4CVMKsLAX/Xfpdijzng33jt0BwA9G4
ztccvrqG7ZZEVJe6+m9JRGvOE/GumLeSBnC//UUaKFXwp46qYxUFt2Yk7K8JdhBwssJzYh5dPPCT
7irKz5wGAh+NONGgwuiy1wVSuluna9vpBMg4KEMOdSzN280TIV7vG5XwYxQAp0Xgzo+qDgqe/Fw8
s1Zyt/9C9BFcb7diPFcLvuUqINV6z7ekI4ZsIPozBCxn6/b6bncbzr5kXv1lEVoB2ikpCca8zFQi
VLSUy3HyGWg6VoSpHaFwpXM9G4yuoQAFKjSFGS/vYIWQzZEdt0ZPG4ulZYc0rbgOjPL7+nfpsHXz
FOTnZHi1O1Gyj3Szhn8Unfjv1RLjQRxcf1mZi73GAv+cKozT9FVYCbILFkxzZnZdnugn+bgKUgTW
CTX6RcX1mDcgYRdlwGYUOKiDzAxlPKo6nbSvgOdjS9L1Eq8RIyP3CmSZKwc+c5ir72N5gdiFKjwc
tNpGzggC4f3QalBQLaxF5xxVefeOrTuhmD/DfKMcYI8SCRGmQG4bVJKd/k9gofZQTOAgrzWPusVt
HtLg0J/Gnxn64Aidvr0Ob6r6ARijDKBl6kFtvkIURRdLwpwQ2RULFkelpdmPmVRcN/fOTiy9yuZM
TDMhHgnWUlZd8MHLW/eKZYIa0tAL67aAb1oQDalEjk6x5ZtQNwI/ibeaAbnwAXYAXStpMuT8pavn
OdIfYU5sHo/abanQLaDC1KX3mWCodaDmabnZM9JhsyAYXabQtO5j+27bfcv4zUzz5U0ssPzqMtfj
00PFVK82nhERQ2k+2GPJi1uSpoGk1J3HGHAhFF1C5qnFg+WU6Ldkryzghc7XI/6xrDPK89hmpESR
5FwecHckDQ9tjwF0lL8RIGEO1+fCHvSI8HlTveY/dbjOHmspqeWdSZydPJlT/ZX6zqW2FG/8+iJP
gHWxP7wLVmY4vMikQnTU9d5rpVI2AkCFw62HQELemosBxFt97O+HbRwl+X97m7nGtB5BeEkAdNhW
VRO0qKOhI6Ll4Q2+e12ZUaxP/gGHuJRcbtroA7wyLjVdRaIaZWFzfoDZ+5jII1EeCvvLu9Ut/8Fe
F/GDd8/YITlxg+d5arPr5uEH6uq1mJrqfceXi77Fo0FUk/x6JizR/xdHm3xqJQd3Hc6lXfeg9dcu
ikAAdZHIglcmfi6p4b4qBGy0j2gIFMNcU6om7+ayFy3RYPVqpFz/3eRk5Fc5QDwbSjOWtR1IoHyN
kL+eLBybZeh+SXjQCEq6xGVz+Y32exlDmwo1t/6h97Aim6MI/VoPv0LeVrQ2YK/LmRQOwJk3y7XE
0sFfcl8wQN+NbygAJcqBbGHBRodzHGEabG2tXZpPEi7KLicFreVbbG5ZKt9rxuE4zC2IqdQkzja4
TpTEgBSYia9U0G6DnmrwTmmwYcp1JOKp+aaUXe//hn7IrfkCAWvzDn0nAR3dD/MHsxQjN7A0OdUU
cue95skxRmIf3XBIim6SwP+oB/UNtizX8RYEHaw56/3MwD8gJut4czt7z/uCDrDpqjMnMsPqZ4U9
PUD8qZE1WJHWsX6JMebruQyiElHapHMNKAsBhUnUgc6ec+x5esShL3aV9sd4XADYqGEpxEq3rdwc
+gb8H8lTPp7s+y6PLqcuhXMYB8HOHmaVsS0m8WPfOjhSbjrITY5P/m7G6cctiHPbAthZVjAExLVu
Ev8AzYDCQe6fbuCIfD0dljwcXCm1//pmj4p4/Jq7FOEysPYLFPBKGEpuzhKWUaUncR5VooAAfi1h
p0GFhnoqvmcUKJhZC5h1UQxqc1sfo0Y2Qni+6KYF2UCb6sOeXC0nh4MmdvN6XUWz/iA+CssjHPIu
RuVfFkQPOG+t1w6zcESzml2/2EqeHlTQLL6m3MzdUXaSyaHaUhAqfItW6UeCaJ00r+oQYzvNvjw4
aJbs50W2xGx0zJ3LL/JFFRmcjMfw943ws/Ip6AmQf4d57cX/GJKSGGIDVUFtIFqzmO9cPS8hxdBT
U8etaArc6RmDDLlIMsxHo2lzCtSFMrRxFYwutuk/a7B94+jAgAOU5HbPvleFL31NvpmCx0b6HFJl
0sxbXkVloI8RJxiiOLjJeMzeb5iZ3gpxW2muvzi2daRKT8M7vNghVGokj5ybyDm+iPoItTfI6c7Z
VAI/DD42mirdkbMaP5bs79Yd9r9CU/Sw11seL7FTIKFamNYcKZoXEWHvuQ8LVmlBSfZg1y0RXDo0
Zr1bSxt8rWDLtCya2WkuXQECmyg8KxMSrnkQk+bv5ceFN1xKe85p5aKk/3Y/6Zd3ypDR1FR3JCZC
1KkQbG4WTtzil572XF6JUJwpy2xCTTbMkPyojZuoWLGQGojs/Xq+x7H2rc1DL+fWLrsAiGwgGWvj
tTUYrkkRShW4rI9Ni+QvJWPEGpUiIROn8kkyLv9LX9EeqLJFtWZQuQY68n+oRu9VGYfWFDUIVjb5
xzqhxxrE+jWg3DlFaT4FnYd14g9OC52RVdLlCH9yBqdMYBIOCzEhwiLYhHI+ht05ZpQHNdwI7Nvo
K48Dibuu+EPmgpmj7j4nvLfoH+IdVkxVLilrY1RAgxmi449rar871LRr0Y7vgSSRgsmFfJpk9gZ0
sx4YbR7LWxW1UDBlCVLmpEJGNRAmCSj1o02w8Uqqr7CbsckjuRGtFud8CcGgZi/sYvTNYOL09A83
D1KUAE/SN75w6TZ+weMkUnW5d38vybi9cBG+y6fGzaH9i+2Nzol7b2NnoGnjkeJA1NdNzC0ofZoE
aanhKYc4FuUIRMc2XHe0fFMldb+akIPbqoB7uEsd4RjtLeUXYxY1M0nsk1Oy9K/2ZaP3RrtNl5So
ncBrjLaZiwr6NeQrBSDAVxr9wTXQwnFk/UESWbiqoPpJqjWTQBEJQQ1fURdldGmDDziOQzfXV46h
fceyI+U2caU+Q08yt+GYNwWzYGVyx5ghzxkgNz5Z7K+H6cH0qwqrzP199GBO80lEi2LC1LWlye/T
wpw9FO1w8+kge6UhuRe42GgIowM3pryrG28qxX0UEgpbPzPnNzmTUZKWavjiYbOYtk5cLng3GHBP
WpH3Q08CuQXpqZmVVC16B/jAo8TS+wWHXbq/7CSb6FEgONAJLKkG2/QaHw1+XXru/oG+JU5zYsCJ
Z2yxa/74mvAnYyS2HcAG53zyDU9NZyIpgVfSBzeJg7VEyW4PJm6sXQzR1tm9u9V65V7ruvumMVUN
kz1h3poRRG5CBsv9ErauGuvRFR8xtNX2OA9KyudtuAoIV33QbMxqdXu2yWGfWZYDkdqWigDsXnzi
hiRFyZNVxhV95FvbIipMvNtM2vGV+aPcwxuJnoEYGTM4VmrL4+HOdKF9xXaCn5+ohciespKjf4yS
kiCeBeQMaJ/FFBhQUAkz0iRXcgpN90yrn7g23B604AVa8wwZwxiwWnLeCv46n8tZbVcGqm4iMdQt
gJPbFNQ6hoRdQ6MrLwUE3Dty5Lqx6uuGVwOe8UEoNGHtucuvrCFnlnqjD5GLb5nMSvomkemcszQI
pnSly7voGfOplOv8SSE+YqtuzG+YwzNkgbSSHBlPCP29SDKaoPRiWRt0URF1PAjVPyyc39a38UOS
mJFz8uo+rrO+FgANH2ZWzhN+4uE0WuBv4GpN7WM2HdP0cBUyAjEu8/khvroADeLT2jRLWnM5oKbd
+zdscDjP7KphUhg5+pjyxxpCMHA69KkUJVhrc3cXhmTIyo/bvOALTLWpUtOurx4i5w8Mu8Ni01hi
TpvJ/ajOfscmR5BjVPhoPnMCU5Sz8dnBI14EsY0pyvn5/Ca3W8tbS0uSoymopQxd1/mQkjRdIKYR
Tn4DQ7QS3UZMYi/J6xmsMJ1S8c5fknB3bSDJDmJTtfyJxTo+ZualhREiwok3CKBuZ7G/ywq8hzhJ
YWWwpZgSSrpro3PSN0LQnGLecSHWp+RCnYzR9WIGDm9ejPx4lPuWgg2Ze+MbSUw2mw1iC5DTFdv7
sKVfbnKzkCxjLPoZIY5NqVVzb1wppJQY1ip9Bhu9LuY2KkI4dW0dU/jnkBs6fKcZYlde3IS5BScL
JjvFOvZl79/CKOa8Ps8uhsA3jVObsv3ZpAhthSDZps/jssZYKP9hfBr7FBfqOLydAB58CX1yCNBl
v2DElZ/N+WYbnpIb6bzR6vlzDxKHfAEnCF93WCjyN0m1gUnhddRdge25Ii/W9LC1ES/cuVVu/pfY
YqgjITSsstzOnea464ORNhbDQiD/BHHGWlPs6ZzcLJxCt2arAsSl397wgUZN2VRyFXY0gYle7Cla
ENcE2fqlywyy3fLt/FXWeye1vFiCkvJpU6NLd3UxL1S4bXn0M5dSn3FryaykVL+rGSdVOxZqugbn
xD0Ksj0n4C3sof4cSWvg6b7fRnDPuSdk2pCu+1muXC8ud4rDW7mqkAFHugxgUeOlj9KpBFEoUAzX
yPsVeEsMZRhF84wzm6UBGnLWSt0/bsInqMqgmjBRItTmiwxOTxMAFJiFWvTS80uYReFkhq/DxvJO
U3TvjTCYNW9tYYxreYCvA93hAwJ5s87PDHpKApNmaCbJVvDyEF/6w1Y8ojznjHn1FrzRQJu6ss12
krHU6+euZkuiiCxG9j3eHStaAwVrP8u+t7IgK8F+Rz3LxVrUK3PVlhwRyRVDamLictjkVmYU/Xuq
OtvzkMeNXaOaRMBrFkUyJK1d2Ek7eeJuRDms5EYppkJtKi53Nyg/CA21cFlQAIpLTf5HRBLDhh7s
tOAznVdtI6g3PuNwtEX/c2OeM8OcUtLEj3ZqK86i1R9EyXcuxnhItY5bG4nJFTs0p7q5vhX+AjXf
zL1HVqz/ch8+bOVhzFQP08UZcU1q20XJAVnf94aUTapNyDgy2DJmyVITKY5pzpUxup7931lw5w9H
cNom+pPaker7tUmbd/j+E2+FyHEXaCYbgz4YXHWt5EricRKJD6UaxNkNlOVFDix37X2AeppnDnXQ
f6C8ViFcg29BHq+bYiXgTUT+3SnvhzEgZxAIOnfkYj32NmV0ZPtouMYXhSYlC8R63EHd0axprpvI
pUEDhr6FF54Sjpp1Rgq+/yJdIPiRQ4tQUQGnMZTqHQjPQhwF5sXil1tua400lgYy0B2XpQN933O8
wp1aq8i3V6C5UHeD3L7pQ0bb01k0G1Q3UpiwutJiEJr8A+AsTuCTRVgOkZVh4lxyvBqzV9m9pwJ5
kxPOd5B3JMfUOoUrfu3+n29hihgObNE+Vkx0YUUE0I7egJoYPkEL8xwh8cj/yiVD6b+y9a5Qs9gu
Cic5NRmGEp/g7u4vGGSj2mlTwZ7yZm3uk5nBbtBRJsAYMPmo33E/7QEcWdASIKGjryiDvpxW5ZdC
VPVEyxaDuowvqZ4yRvjr8BxwlRH/eNkjddmnUGKWRcDPqqxPsOAZ1NNvwXsHtbNc69KtrW6MN0NG
RGZSGhrb3TTU2z22qLMIL28eZP2ANvc6AsOpSi1HkHTmQdU2DZIQkLFBmFXRoXGxSk+LYTNtz6d/
YIeWYzScXY/qlEHEHknpwKxswa1S2l/bzUEa/8/fx3VlunUlnM2Nc4JT7n7uPLApNjbfQ0V6HtAL
BSlPabuNM4OLFgPSZ3CjzZXVg+XG1CSfnSWOzf4KlUBAMbb8vpz6PqB037yfjJiVcmp0pYyYpveI
Mce3tnsZ4455P3XPniVmhZ18F+v20cghWZgufwNLiO0DRF0TPJ6JZGK6ts0/Q78utgx8BysSvOeI
omNxa1pFdCnMjC8Z4J0NUzGnBx7KgVVgVCTbQGyKqy90EjL2Nt8bAtOLPe26xzBMbO183wdUcoSF
xDlRNuO6xHW6h3014QJFWF0HTYcU6k9wQWtTjED3pUTwlhiZW3A5RaY5bRZLtM3Q3ol9lA8xnGQS
qW+xCOWDRtR+EpjRVVHsPpAgCgIatF2qYyBFZFuL2FUWf3DLUZW6frkbHAXI/hh0AyCa6I6+2krH
i6RdJuKjbM7B384TstJffX5N4mhgeLroEzSPEMzqa0u8tIYx0oIXMrsm/AXfHxN2xVOFaZcMqP/t
Mw+hcoupkCkm0OT1iWFzM6KOoQ4OgCJhGow3bjvHvEbpbQ1lZaYP32XqnumRPZjCcBdBJTm9grhT
nKQZ/dUZ6UYd2WXTrUD48zQwYnUZSUJuQGfC2da0rtyw/q3L4VeZBIkXnhQ6sZ3JWEUK8YaFL2aa
7rNR6LjZczRUpQ2O5jOfTS4kmg0dw2G5y6Vas/f5AseUxZB6fHpyVNSsee3UTPEVQdJHHDLEzuh+
EgdrFxSJSP+2SwoveJaLXQmrlwWf2zB+njtwSeDE+z85ev9D1JzcgRhnrKYCt4N1YxaVA3Gsu6pS
IxSRVorGXLRP7E4Qix/0TdrG22SeLhjvIwTxJbHuQtfB82Sf0Ycm84lfrGnwzt/SergCQhW8jejW
AvNtLZb2q9UWcOw8PZ6IxThJ2mdnmlEMfW2SGg0sAnu71hpMeXtb3AEmnmQFVW7/TbUIjRIOdRaf
yz5KgXf3JZ1sy71V7A/bdLjb8ceCXFKflj8VDc6XVCxjh3tR8/BqXjV7uuJQvm/pT3oYYl9k4CxI
3HTTDoGeU7y5gLx6HHfc0YP8Q11UrGhvU3XvxDZeaBNY3PlwB9NSwd7Go6qiI7ZtEJvHYLWbdkcm
wmxrpj/4y0X0MPJaTEDDXX78Jcp/KV3WPISty6VB5TT6oQtdmjRPvPKN74IcvY6UJ14g0TT8ntrM
U82F9Nmaduw8EUZ6yZPb53Qv5MYE1gO+fzK9WrEe1RRDgOd39GOeWGjFLvylpbRtSUsYOD/AlKXO
Q20Wse7RzLUDQ9cSN2/XlCfY2iP06pRYISmppj2dJMTiSRxfSLX+PRaesADqinOu4KubGXVrprX+
YMRX/xAD8i1ytSO0IkecgxfGeQhPMo9JUv0LDFWL+Mncwsa0C8x3BEWQdxwH/DvETnucTQDDZxo8
NmQMt/2oyU1gpF6zQDZqjjiVBIJGm2UGiP74sxi9sOAtqo9Pa3E9tzYWC6+D5jdpuZVYpr9b2DSH
0EudIcKWy8QTlSzKk1SjXSu0BD4/bCqh+c+2oBMVAvSFCuW/a8ga6BOuuqCaS8SPfTVTnuZhDgcm
OQKk3ZkVY5F9KqNvferzqGdSugsAeY0yo3SZfBSSHaXTaDTsnzSKhiy09n9USeGDSZJGhpWVz7f5
mvnVXdvUZJ/Ia0XS3Cp6su/UP9jXi1nupGpzCSQWq0ALhMXTatdDmqtT6uoofzR3EQbY+rrffp8d
KyDUG7R8y65yDvTHSSN0ik2DyDKVAIbpkrSLltflWhHgTUitO7Pf6+Rvll1PL2XXzd1NXAZrwhY6
bxYZJttaJMT3JO/GbcRzzmswt8ZXJVTfuKhFf/Rhk8yPYQ7iAdkJVixrDepiSTtjslq16T6fR4mH
bYQ2UaMGHPpC55/04hEAhWEqFPwsw27pGZWK+oK/O/TxRviSyRRzD57IEkk1vrmhMdy52UQyO3cJ
AsC0UfmbTdOoLZV6AnBx2Uuts9VqzUKRaNP0q7AMrjf8fyLrriMopqBOViJkbTHC5j9WeK4+wttA
9nuuf9F5QDkxP6UGObWUAl0otB5K9XK/Cwk265EGXP4a+m48kNQfaO/xnkxaGS8/yMOts1jKJNkX
uYR50WMsdBDSRA4CCumVEIzrBVf4sF4vfh5A+Lp43dhPUrS1CNoDy7sFjedbpmYxyEzc0HArSiik
W3vUHvkrCaRnHOqHh+hE+IkBZ1Rno08jfNvfPShzyH8YwXdZyroMtDMqLxQSZE7FFAvgP8UB8WMB
mCUWTLBMOLZf4Taohniy5K9iLVWSfoxkR5WNLgxBZg9rA9529gVAWy32nbtMzqZXDOH5DanEP2WT
q2keNvpD2EwPPrvoNxPMpy0CH/c2Gp0eJDIbbxmuT9x+Y0mHFmjIIdqZdt9OFkDp5DPOOtADydn3
ucvbcKxFHZXxO9AfrCqXAeh/MWDgoJ4kbRyqMWdPfK1uuZCfQKNTDV42o+HwNXh7CwgllfP99a02
fPibrHgTZBp3D8FWNaX2RLSYjV4chWp4a4NUGw5WKgwinegXq8QN4mPi0whFeXtaXK3WEyMiE5lT
SZca6gL+X6czNWJMQkeGOOdas5QUpNuEZ639toac15fbqt78c8q26XuFwptXy1CFA6QNCcmN6z9v
ejWwb8/a6lqlnfKmZ4/BguaijBwzEVNnLEBwtfPY44tbvvF8KDojgp9shDaDJQSuSabXvJWsAcTU
9KGnYudIrL+Ue/eo1VADzZ4O8/WcfDBMpPMrWH5A3sMgbIrKoNbhf+a8jaBzqiEELfJ1GC6P1dEk
0AeMWnGI9pigsqkkbkm05eO/CwXUk2ZbqORiqkcz+wJm59ZJ+A1dJfIlUyiPFuovrsbG9U3Fz6Ku
TZNlpPQX7ihu+0oJBbHv4xO2alCFcQFYN6pEqpw4qEJCzc2n4dAwiL0xLNbJOV8nIOAD9hTeyylZ
5AOUaEjqeZjI5y/xAvW3ifWxLyedXfCSXdY6hpz01xNoco3qYlbQtyECbGfJjBCguCgZTK3WfVhr
gq1FkXRlr3cXnoUNuS4zqJWUdlnM0f5NRlSKSGf4d3rWLVOo3BEPxCx/EwKWRiFBLSeg5o+3I3bO
4t4EgOglylC3PHprf3jSFcS+TXIYFSCGFVXje9NXbhDBKpDRge7qHisG2OGBToHZYH+9VCTSANFa
45Zgrbonu7UuqBa1ZGQqAnjsMotneqGKxDF+07EzE0fGRe+N6WilPLMOp3C+6grPrDxX8cJ1Qr28
1l+5Z6QxJs6fj5vlw8+EdQ7K9cHWzzBNa9XZgh74+CkGa+JPKNIYu5aEQXLJqCzYp1Yi9sbHFuem
yuf4Fq4zEGYULa53W9JWZ0NiisgSQ6s7gmOETBgf1Yd1oED8rJiNeJJbZ2Tfcd7FjmzAYvP1hOO6
a2K3EWcwJRzEg9o3HlNX2F3hvinCnbn3PmsHvQqhtcRQ5OEs1mCqcC5z53lFpAjJdPv5vc0zjvBI
rAtqPya4xWX5RwYAcz67pGG1k3zI8JXTBFHFbG8E4oWWasay904E/WWxhu7HPaqt50B2GJq5udd1
c25FFSF67KC0D/5/fLh8eb+tp0vTO1sSRSXXCIGzOj+GcIweUdTyLLDKmoOfmm4saCBmz3m+5Lfh
GryDP4Hd2Vn0uUrEjduLYU2JYe5zlAs2FWwJUT6m5yt1c9TJ6r3K/HmxMgvdA9JHr+ZqDYWb0kj/
tFlalk0xB+1e39xtpjyqdoqqqvBPLg8Sdnmbi3P6Dlqg6tMFy+c14KmkinXiC8Qhznzc5jzyxGwn
itxXakMDkKq9/U65v3UIl+BTgm0Y00Ncyyu/nYHK3rv2k5IXFal2xXkhqZBSiMmWHUklBlMCI+wn
j+1zhaaxlxgnNbpnlk96jxdjbFffQwKiasUc/bDioh4ilYOJjDSayv8Gqhq3eV7SILC+r3bG3VAa
Jqw/1v5knF8pWMVFgeR7vidgoIArcBlzTFl11SLVBVSug1+YtieO7FUilsTkfqTXn64RJTz2Bngk
WgEMPIXO6mJICIq6xXe9ahhpKMx8YVnYjq3e035YfIuNkVFs5SRezF8EBfw6gwPca0FTULuIUfmG
9opYwdPkfx9oE6P5xSbvbRt0Bl9BToRczMoJPy5UNyKEc4MtKpdQoXRRtcWH5kr6eyp44uOIS8Po
t2JVQ9ml/aXSqcMep/LuOXzJcMP0FQ25ap9t32dx14GX7q0lNv5cHFbCxL+jvYgCrQsdYMu1aIoI
H0dJV9NPbCurgigL5ZKJxB6ywiW3/wbMDyX59Y8P58XM7dLcQJsZzR+1IIfKvZhX8OIBNgN4lXf/
0cMg+2enNJlAgSN+2+Q1+8cuaXly75MO2fDIrEpDIIFrOzqz48xosQegitByNioMRuFIhHB97Vda
O49TNuF02ZF7jpG61MN+zxFqJ2hQJx+5P1jtGAql2aae/rtsEYJnBGFypBtJaP0X+j51RSENWF1S
TjSM04xMow4Z/zIcHW8W70kv1bDkSFq7JJvyIcjnvR6ZKxm2iMYYBnZ6Mq10FHqZzy5zhK/3+XAD
MK6EOYtr2ps5Q/ubmQI5NDf0sDnRYN95dAvAq38Pm6Npo6XeIgrhYZr1aTcNKZZYX4I50tKXUFg5
/EwaeE6m+lEFqHkAMDifrZuPWHfcYJgTbTKJi9XL64CTJk9SOISiPBehWavTrsqReIfUZknPE0zO
GvSvBk6phLLmIRaZHZf/mEeq+VxiiET8uKTtvPx2J+7+WYGr7Skjiqyoi+DoUKDtkY0yU8DxsZDw
P63eeTxt5eet+ffPwdIBB6n/IWyYH2+V9zc3KP/KiuIQoF9cZED+LK/gweTRBjFXvxixlFMIrBop
hAeA3sVV48I9bhvG2ouqNTdfjA3bJ6yTObvIG0RkinhRlUBC8Vt2rVe7amSv7f7KM0u2Ta27YrEC
tDvuoHXhnOd/uC/Hh4cFR2e7FAvoxZjOKZhWtQkXxZQUM3ajSIbzzsfFttERvU8MgY+qNloiWHNn
ojytM6CsoiiVrqaHh4J+wbWijFce4k09jzwnSCRNw5V7QKWzUx458f+I6W6U4NjoMBtE028Uxz80
vSVs9EUuNUDH9wYEF3IOqJIxVHbC028S+B9j6nNcXmWFxbcb9Pt1sizLAfGKZIPntILg0f2Jb6+C
GeOSoSu4o5ixy3idISZeE41VP+dvFoieKolWmEyWp/07a+53uQMbIu4ypTlJXWGV/uoASwI18hMH
gpDwphYrzsVI2rr2skg5T6F95sXBVGC7PvgHpqBQd3qIrftt8cJMdbThfg6BzkSlBiJiwZb1J/Lq
MIB7D6/L6+wzW2iruXpF1s91B0bDAgkJpP1aRvSBx8cGCX/Ym94ZKRtdsaR/v1K1XXfTHV7dIo++
B3LpbJ3I+QNHbi45P69Q0tx9oaI+U224XTwHMztcv3vHfB6YSbfMsx5N8qr+kTy6nnPIOURdfkgS
Bw7WK0oXXXArt9R++AmgzoYxVUVWJpVzdXcB2H3KIYbpRPXOYX4id0sLaGepWRJ/Sd4ZXsi98JxT
hW0Wb1y+/A+kD/e61rN3WCcX6rrE68mNIJJEc3cPXSq4tEhbKF+I8uYVg6x7RA5sft5DNfaRFYBG
omkqyU+2hBZCOnR5t7v7p2kchepZdIAweqqlj5hY4t/HbSK0UM5f0zf0s4CK8mS/Ig1dEQyQ0QS/
IEUhgVTzJ45TMc6BOK3ckjg/0IELf9JajgPHiqknxaMkvDzWCTlVWUmxGO8/EmGmUsVK0y61aRa2
c7QP8vEcW2rxvw5+XhT5/I7mbqbIiVwEeiwMfpdTZgFgb6SCltOU4NBNc8CTvOci4Xu3K99o45JR
2/urn9tPiUnFN9MbX/jg6U7YfpjbNWemGUskA5VEWuHwnqe9D2GNeuecJ/xRNOAqCVOE1GvYnb/4
FjqplTqJ31McC34JC5QEokv4aGO26350BHNvtISsws0jFYWvLDCOSkjuhHEaWWamuSOSKI9D4iqr
Bm2fOK0uN2zEf2I1yXVWcqkUPi+nFizcgZl9atFPWTAl++vX7Cct1POw4SGTFIXa3kKCOWplMRXG
ukfrF9YUDw1wfhldMf3dZ/LsZ0Bh6MriDIz2V5nU9IIEaEf92YkIP8nuoxRfFpd3GsaQpttpNqvq
2uunYJyPLKZJxPSjXwSoWVavNcxmAAbKfpUFo2hFGmUop//RN0Qb6D3ccicLATWf9qMs1xe+Yc/J
5mtulv4lQikxPxUuI9ZpV1Y8FyGYn46Zl6zCoDtxBE1kcSvwTPgCAyu/IfrBGgxIx3KUrj6tmLZk
3FPL3x2FR52Qnos4MJftfuSTYnTkfzfuTRQ7spHcJ1m2rENk9hV/4dCQyzaZCcWYKqxXQokNzPfw
hqTKNhOAW4xYoS/NmeGGhsLV40+ovMfHuxb89o+9SK1Xv2ex0iceDsm4F9dw7nPbHfRbtmZfaOqI
EjzC0TdOGdeGAx9qheeBHDD8GkMLFhZksqWkb21EQft/2jUr+sWNySz7oYgqOwdeCL5RLPJ3cESp
nkzxlc+CZHhaaeqWR0JGzx+hLYjQ1pZlwKvYbeC9aH4GkB5Lg1WHaD0lghdIxt0QQ36uRPDReWJJ
eIIXEmlL670Hwgnb7UPXQO+jiq4EymiPHeow6ojEcPpfxVIrAWnxG7STVzPimu3bSKoivuOb4vOK
AzA+X0ZrrHIznO6ip5okBq7BwnrbVRAecla2jgBvlI93/m8tCSuZC0kbmT8NOQT3nh8XXGb3oH/c
pHdgBu8ZNoYxDveZ9n4+uxZBmbTUemq2jGipdWAqzIkTFjpZUV7glsNDqpUqcmTfC+s4LLFNj/4y
HaThjw7zdVTJv+OIWkbGcQqN4JYRCDvgjYnUjUR4GRprioBrMna4r7nmdX7flKjBrgW7f3ACcUfI
6do087syZ3R9yPPd1pHzfkOe3j+s8z+RQJstSdVq1VX8Lkudf9eUonYHqz+3G2BuFHV2dQkrzbF+
1IUGFaGx4s9JHEva3F21pVp8k/nrakiMN+wjAxcrocMZcj+bGWAdIPD1O497qeBzwRaOiiPVlz8e
CnCN4XtGKtrCx8J7ztJOY5iRq90871XZlTIXcTJ65z9CZJJOPIEtLjP/NuXHg2/HdwbOP2tp9Y+N
AF+utrKZ1GYrJkeuvNvSCRALPNo9uCbv8U2rtbo1DV1WPRx4w1xrX3WP+iz9Iiwoe4zBTIIL4cof
mkaj9+Qpmzzlw31WoeGHTdeRg79hv16n0Dihzy+Vo66GDybshGfnW40i72tNBKgGKcgioBwcdBlT
+JJEzpeCGNUwd6DTTp1plj+y4QUDraM/5Vc43+vkPbnkqISfxmeXyWGJ8xIKIZXrRG83YbEFCpkU
ENaJIGbUqMDNe+IbhPlAtnnfSZSSYSuP3dJU8FAoB/9+3QYNvS7jdELgzjQcWI6tfJOKha6Fk1Ia
YqMBSwxbFtXXal7vjfbZ+9fZjQPBne8og1A3kKC5VKDnUBy17lV7a0wCDwSCLwXgQvB+jYIT9FzW
GZC2dKs3FwWQ8IyT3TV5HTbm39o6tL+bmqo831Ox+ux1RHwfMH5VRHFXLX109sUWmjPYaQdsR8zk
cUWna/3u8SXkHQbXoBjwEOF9tukUCWs4+uzmyCKnxeEoLshowxh25wb0SSbfRb+0N9n97VBvpS9O
mT6+ebcLfSMpkAx85iDtttp/eBffGHR3bou2sgcyoR0EP9Bs3d5LEsk2aDKkuiuHIzVSGmCOOvXC
Y8p16m2QKFN1V+2Di/eEYcWs3SNu4sgO6RhL1Mw4tHuWPpvWNlFPD9JZM14+ljfvj3Ts0rUSXMrJ
bZR8jA3lwSUvqRG/AJlTEIskgGnXy81JrOUuJ4S0ytsvucNGoT/v5qqhKYLG4I+shOuSoG+6vggS
CMNQaBnu4WHThoIDWX4IWKMp2ChQWs/eqDH+afYV5ikLxfXxdFZ4YLqd28yqNQJpoAzYTL3fgM/6
AxB+DOqPWq1BAy7SnPsR8p2fuJ9ZqFzljEkSzdkAL34izc5pBShp+MK1RkvP8gwiXLxWSoVZPS83
wo9mA8QAl+zU1KSFwT4ErUBIx4rBQyw+ip6fb0lRHoySj9D28U9AnjnIaeR4T3xcVkeRaBTh/xZE
tFYVk0/nyb1zKAiq+2CmuLTSJzJriWBtTmz0LJ6SlqlKTQqefwIe1TexadfmXrZZDddNZxqQQHSi
XU4D0UxG3rWMSRmbNSMJZUvN4iMNgAR1WPDImON8L7PfN7sIrDU520qwfta0Gk6HZxAhKgbA1TrV
fmPEgxKu0xqi+GZi0fV8z25a7SZTieZZV/HbYzWRadJn5sAg2aGgUFigTUsQQCwBQYKlSKiOp9S0
vfq3t+Gi+zpBQsf6u+AKkd1UYhI1g1ImwHHUxMTgQ0CvTnpBUzX5SEU0D1UFsLqK7d1Ae0RwVIUL
lqRhd+yyV833XdXVvmBYXs5u83K4Wy1ZszN7Y2ygciM7QNCjL0RnmTFStxemm2DYcDpvV3HPATKW
gLhxQ2419o+0esDxqKOLp0BJ6UwE42vojr0+DfOTR0IoYY0HLWSLfGEHZLNJkhI0AG3HTgErEeRI
5HGgQsXYYIfrpstPu3ecvVdqqvKfmVK6Ca9mb8mFBt9SwFaixeGJKoO7P/y8t39MzNdspNwcqfPM
OPbicn6oPjbxLYt92BZVw30L/G9shmkkM55IZdX5klNCdYDCO2xFCUXvl4xMsh+1QSdjJvok7iTp
Bu3VgU/+dcBjHezjrHSRp9wjIQ1GtDDIp9UZpnZ3l9CGvcaOkwEREskOC7HXc8tCN3+5FT0bVOrf
fsYL8Jmrd/sSvqMBED+9iBAL9FBOjBoJnLshmYJqpB4bjHPqXEfaENy5qk3tiF/RZZkCUW2Z9VQT
y1UDC7t3LYAmoM7kk5D7lletZGLUOFS+NftQ0jxtzcstPj0JQNLiMlI14SPaayF4d3Haaf7y4GXD
IDrHvKFcIFyjLcBeQnxbFJQUJIKjvihAq1QEexzaNS0lk3mkdaTvvaCRnbfP+KaAFpNr0yaVUBKr
FdescF5peJ8+nC9/Sq766QmhftiqLIIyaf3LrQKgNLq4UynAWJQkfoh/h9fa8mLM+vsrfZzGgz5B
vSNC98r9uSHFzKrtGXiW4xv/RxvorL9f7WyrwELwrci4wUcPwnGlFfyy7NGwwRbnAZmBgLYFAry4
N9juoL77Nm0Vv0cCyRSEY2+bP4YbsCqTHBXads+k6QNazQRaAQkkGOOgy0szWvvsNx1maeoKom1J
4AT0fkgdlfTwuZaoksD8PeN6V4mtAoDAXdFN/gI564Gg/dN2vpzH8scrDm6hziU9BeAiC2D5ZS7+
/UrtvZMa235tQJnDPVUw3miDkZ+z0opVf6QHdcQg7gBqDywn9/7sLQx0QHDUTL31FN+gUn6tTp9J
XTQkYI9dUrS0bNsy58vZAIvbtIGNWw/Zkux2maCZN5DUWs3+p4NXeUTwuR2MQS+7gPc8K3YNh7Av
81cGBVq462kzFr5vzbr/uBOBUvMoBVHksvOftZ4KJcTjTUiGPXQbhhzgAaszRQTmiKdc3Eg+VJCk
bPUa3RkYxMUTcQgc/lGO0i7+9+vRH0Ef0yY5qzPwPhZI81qFdl0lYV6D24voO1XpI7XZ96V7hWjt
O7Om0MR7NHjrRNos1VaqXs+xZe910NcR5wwKTHQmNr8N3D6HfIwA6Ljbm46IB+9UgKxrBT0LI5u9
ulpygvOvacJPnWTU4PcDk3NXZt82n7UaW99zDkSNg4clFDbUzGrqQfRXlr3A0mYxVg5iCgjHd13L
A0u/9/QCQvU0JDAYCj81mHyhgLyPD7vLnGUGJyax4Hp7meiFY9OfFDhR9FECqq0PxJX1F2sDvhy1
sORCtNgv98OOu4OQEKDmaUUN+PJ6C35YlYCNV3267gUNN4/3VIJEu9+tt2n7dFJLWHGaFBvDuZWs
X0dVfXvMKlFIpdEfsCjICvg9yOk4Ar3fe7njfsHZO/z8mipyWLh9AZHop2fn1h2VOe6uX7+H2WLS
U/8uu+Yqz5hu0qnEfnPzLtVLKVsIn2tRfj7K6+9LIUdNwm9OEDXkCVHNFEwRZaKZ5J+WBMOZ10m5
/+//LwrDrHlPqovh45+9/5N11syp8wz7BA+Kthi6eyEHuGnNG26rODmN/PJ9VPyU8A434CwRs7/1
GHAjEg3PE3CuVPvZD+hXvRqsr/nOLkUFXjbaaZoF/N2BIpsr2IsaWXZqwkev1jtuCuPOhJ9aHOdN
ceFGzp2WT4aY8Lc39HtJ7BdGducFjxawnfxYwzLkmamjOEwyfYiQBO1wFzp8je4WdB0U97aUnZXR
XoAcFujrvkzr1+dNNfoPbnxqb9t9ZE3HCvMbkQJKFK2yERIJTzURny015JukLyAT/aplTsRKbAtH
xiwJuJ8YwCF3him/N0SJPwNxoMcAFlDQG5HzmwuAi8ad+15fRHKJ3+zihVm653TUo62gu8/B/aSI
1wf3s0y7n/L6sQnDa/P+YY4mKsJDV6wavcEg0VJaLGBLgsnSayFCAQfMz4PM7GYAaGoQdaSvn3p0
0M90d0xfjGverH7oJoyVTM9+R6ohDlUT6M+4yy3eQgOCC7WNlZj6/ZpU/UAVzbMdV9zT2zPUq0k9
U9SeRwWEfKEkXJw1+/UR9WKOZYV6waRUc93IZdb6eEA7SD5s67F2bNj7vQQpJ/hZaXau6a2U4KfI
34thSPuXjADaKA4ttVNEqHT24MkYUoyRKlTzfTJdR6C5hWLz/rNthIOtabc9rTAtzRlORJXgsgPp
uP1y4LZ24OoePshGltA7l8/fKvkVWHafomZWVO3cXenHwkAnGzosvrV3nZR//HunIhTudrzvj5Ed
POkA97c1rVvaA+xMgDzIcKQjAwtxgCoQJBWvkoYPDqJP8Wyyg/Vx8hYjLyEuvzeU7rGSH8/iCVLy
WVbnxSIc8aWgrwkWGkobU6ESK0ALph5P11bGceJ+5iLdUCXtyuc1ypkjOJ1A3hvRiscAgtwQTmKe
jiQNsSKe/UY7hgWHPIUBZrCriw9kjoV0eukcUh75/FDfVDImlBeY6XWL8uKRcuk7xkMnLbaOY4ix
sFbPLuliPJNqCSAbsUQdPG2uzr0zaL23Nti+Z02NlrOFx1kwGymqWdEbvoaufT4wtY11UBA7ZLoy
CttIVoLVawizcEJOC8sB1hofqVvlUt1GxmL7BOfU0TKm/x3CFSHVmpCgWlkjujFpx5ZHu5wXN97C
hOXnDU6OhQDvc12pJTdIgYgUpxEBvVIuiyRdXp4TLHhIXZaPNtrMvXHus9isExFITjIgWCDzbnsd
KIuzdyZE/U1RjxO4YsfQxBybpKrnvtdhSaSOWXP2EX5a2NzJBEmWSHyrB+8+yJn5zICcmkvMSXUE
ciZVjtYJa8OAD7tAw3H5JDRUG72YxKdgL6q3EkfY8qNcRbkG4KLnLXMmQizJmpW+n1DNhsOUNNh6
d4cRei5K1N2OxQZelemdc3fWJnAh6rjsq6gqQF8/ePWH0e5UTDeRMrNMxp+v0H9bh8zB/fI1NNMz
gq4yAbPXjOcnDuVzXK7bDzS1tLJA2Dr/iHpAqCwdL3nMH8S3AI4Lq1QVEyHqxDftYI1lAu8MudV+
hmbdpuFbYQNdVPS01M5P73OfO/jxD5T2oyoXda8N8cSUhovaZEDUBJh2kfUPrMcb9yfPvf4/qkdz
nAv+GLV3C6u/ytq9cXzuK4gMKtb/Ynh4Lj/AnVyvG4W1/u1KxZbXrt7WUWx5G9w5Q6RVKu37T/NL
wXwJ+T+km4rXiJK30qP4z6h36Y5SwGz2NFLaTujWcGzJOk8kNrDp1gDiYeWpqQH4DUMWs8NeVq3P
ZJfZ3XKMSvuonmEP+UAan5QTHok6oB4UOQwxZWUG9I+QYVPx62LYarcvxeiWpXtW+63d8Ax5AfuV
DrLc3ggUv7kfGGxeehAZquhzf+kb2APvM6962oN881q0ulDlYtjINXD51xkCzAc8ptjtPh5cYsqC
iXdTxDuzCKEm4eMmn4DPCa2DUgMSzGWSn4uja7Stiee6xtRlEyLt91oWEUc4vdZNyyVv2PX/TFXG
4K3BQpa/u6t8b79u10/W3Jhu5A1RqIha8+8VB/voJWXlGf+e6Ggcb0cTbpkGeGyOMh0Ww8wjYVkP
rAfyIhKaPmbcsPJkaodgJMGqacmWNvTQQ7yiFfXI/PQRBF7eqzfV3R+TVhuZvKaM8IVbseckGOtU
opiLDBq+UBNVFcdRIIwx0xSrAQEDjeeWRBZ3zU6kctKKdydsup2j67poDX8F4+iWxlVX6urzrxuj
fH74Tr4AbLwXUmHe8M5n/726tFM6D9IlgoWMn2yJG5kbaU7/WAaB1z1bU190egEhdauu4S/G34ug
fRFpxJj5/JccaRHVe911vqk6WqbQr084dU/pqD8tfbX0q6IkShv4a7tl0HuGonjBYgL/QUTWnLfy
7QlXrcBT3r29uLhml3zmEfAh7EnGmEEVhRcpGs0zWp7K1aVVl4YWMuAjqWztRySqNFyN9vgMYWRx
yAK2CZHf9eM8kq5Vjt8SUG27RU8rd1S7gmuYp8/TxRdiDb/e2IKHem2PxeXfKaok0CK+3tL3M//+
tu2CbslXjAEiU7Zux2rYgctEbfGbKYXCZ1ZMdwA448pIOfddQDGY5YYNOG0Ch+o7eJ6AQFcQ15ep
srCjWdnQdeteSzTRvzFZA1Dpr2EvLURO6SbgCuNanG/84QR4mH4rnT+GezjTEdcP0K+drZOJbSBh
6UyaQHCV8JOpHO/7EaGTyfSpGshk83O7bpvYOZ0qQxvMY8lYem1P1dfZOb/P22YIEjq1NxpD/zrU
TVlU9R8RFb2+j8mZHd6HY7JZSetQRU79ebnKmHxTX08XhZtC4RDUE/gJG0s+oqzK5Gd6sgLvgM4H
LaqoDon35HNqDXjOHoPvR8yvdk3Ymyx8jikwskZt30lSeDqmgXNYYa7mB6yL3dTswJQvZpQAir6p
xPV+TFK3TdO6HSYlO0nrRCrsXp8qpYXtxXRK6pFidWyZPJEFew8KzsG+KJWno4s3RNFoFgkhw8Zy
Bfi5soLjahb6P/4ONzgBEjzFdqCDIg7cKSIP1tqUhOvl9uom6pA76NyVtAz7XtdZGSEmbyYCONVo
vTGpFkCqED5UB+Bf+U9NnBqraZHaEFvGKURwdSuM2oPwxApPqreNk+qOr3Twyt9zH4CLda1hHK/H
GvMWY47O3FtPiu4T5qZWkti2+/d1ZW0dnaNKlLH3fqbjBxuUSnKXLlxgg/+3bhYCQTUQVHT5Piig
zNYtKhjSpLIgA+UBYepyqapg5WOsow26lEDVxi6wcuUROwobD7Nx+NqzxR/2lFVl1i1hsrBW4IRR
AIgBvFgiRjOde9rpV8ubPtR/TCYuTij24zkPYYdgJ/qHsROTgcOH6BjxcKKyY10SXghRkEN0DO7K
CV6YY5yknizkpHY8aNV22vj7SPmaE24NzLLNkxsBB5iqRQtB1bf9a4qP8Kmqs+4ICGkh+6Y9zkTA
OOsZIw/LnJWrT6bbpV787jkq9Jhs34gU041bu8hku+Q25fI2zNOu6POWMULbaOy/N/6E7U5shaUW
FcUrwtoRuU/UR3hpTNsWhycQkq5e9iN3iMx6M2Yp04mj+UFRJKQccA6/jhX6jRvBpL2Gtw072OQr
LF6ExmYe/d0VdJgXVY+Nr2XrnsIss5a6k7f9Zs5HAqNopofFCLe4njVXa6WtuIUAlwai0aS4SCDU
b2qTSiqTvhncAzUUGzzYWWRSGPVWmCQESXF3ilfiAUybCvgQfnA0zDt6N1yAiM09KxR4OTCeeLga
4+P7YIlRsSyVnZZYY64E9l/Eh5uJBkpY5dLLCiI1IZ/GZY2YhzeXeMUy3VFBHiGjctKE+a2sE9ku
6K3qiYVDxYzyWOm0hi6xLKBZ1wgYpGvcx9h8VdRFlY99D1qOO8b2WigXTXgMCNaTusOLDs+NjrzQ
LkmvM1DlbbMkH8AWUKZacko5ajt1hGzzBUwBf6XrzUaKjb5L801BMbH493Lrl6TgYhNqxOJCUjaN
QSo8XTk6hDtZeNDglPCsr4i7o9hvyIv9D3LGlPC8yKX8NRN3xokRd5gKY3z5i8nr9rZHN95JkBAX
EDnzfOKIBoAbXdAU6YhiVvQVpoYmMb6kfp2iS5wB+0JMAjVpZuRP0A39nz7pyW9F8sJEDATEpfpo
ZCe17Txe4YEP4/6Gx3cLGxOr+TGV4zwzvH9DjA88K5W1dQXv8bgDURgGOEdgoSldyVm3NmC17D9Y
YXw4MCNrLNc7P83aL3YIS9Pmd8JcMy0bLLHdHtUN5ZePkekbHSjq0h7kpsuh5JGoCJDoMw2v/qXy
URUgeJOV9BwlssT6B5+Tfh4bnQ6w4BalCTt3uSgST1Knq5wfdBVCQpQAnrZakJvyjvZMV/4dPRyS
TDSyLLh+l4kI0pQHG3KteQB317X6DOplB11imT8TV93/dp1jiZ5XgxapivrlDI/VCOtycUaSUEY+
YvgZQP+rYTy6A2xiaRwr9Y7gbchTaNW/wXdyUBCn5OwigxcDRIIwLyc/E+dM5J2wxUnVPRDWB+w5
EbFQU6loOopMQLtvPuMVUbl/mI+24ZX9X3A01xY0E4+FCI7/DVoqVtWk4EpyjmVfu6iEwmUAhgWD
LR0uRRh/QXHcV80CIbrij7ewY1QwFz9JBR73FCkUKXGXEUe0W5feihag0z3RRVwaDlF7Y9EfLB4v
uxAS21y7IM91doYIzXDk9bHpuR/y2oO/xxYEuYM7KV5Qe1Fz+rc0BiDo0efdkDZySUSvwR37Bge6
NViArytjMFQ7Yykqd2eA/KefOdPZc7A5GePikyo4ZjaM4N1xE2ogwKKSlDg38U061jhKQcXGsof8
2ni/a75y6h+O1FQ1Q7ZNfHtAqNDpXRFZ7UjkxroQW4it6TkeICT29ngT/qRtu59fSIjaZBoHiDiz
pUnG3BlJ6BIVRJ1Uh9KWDOtlUtF1zij7j/M3bOT8kwd3VJ3GngPY1PMqcI+RW6CrOLlAFXWUxmE5
T4DN642DpSCIfEp+LVAzK9dyU6D1+fjW8Co6aPHCY8zaiLBKNhNS/0Y6wzLE3fr9naxu+rR+iQ1v
JNOCf5asI2UBt7T2K/M9ukDm3YHbbnvhfEuXJN9FymhtxO923upHelg+jInJaQ6a8HgihiyZVsvB
1jowuufvOjUEHF/bYjRyCqIVJ0bk8JbBrd7ziJixFNYXEzOGjXzOEcMfDXw7gypql2pbbA7V5OMl
BJ0XbUVMU0FvryPhtReQ41Ug+xevnJeFE5s+RC9Otp+5HtcR6aZfyqnFHe0hEo1x0TIxIc9Tw/1S
Ke04+5NdXPyNjIRZhchmyx0GksoW7LYQuD2VUzOueMz/gYeX9bV72swgAEiI8Kl6bAbQSRQbx2zN
RUumfM3Fs1G9ra/Dgo2+qT4Lej0BaKvTgmmB6Iu5WN89dXLcbXar8hJDgKQdgIrGakx7BO9C0Tge
msFVJtQmBwmj70YJIhyELVz8HnlZMkJUmasQ4qB3JbnZHv81F8fyaemGIxhFd7iS8V7Mh5TkMM3U
TwBPthbwC8iYA7rAEghU1aiQkwXhCPNGdDPJzWpfrdlFVXt/Rt6f7JmiS0G3RCUr9VWxoYKrsyZ9
JCPaP0xkfmhgxAI2GNNvA/nSF0XDdUwQSGJLhKFEwdR9TwzGd3+Z8jfBsBYC67ZJoXRkysvhCXU5
H0WOrglUXmG9eABRrjGTe4AI6MqnnI5vTYIVOfXt8RHK5Rs52qlp+fP6UpypvRyizhhc6mx1DJVC
7GekMc9Y6ff5odV56ZwZJFvz3n/dBhjJ/jAfUkfHLFxdzLVMP6076Ripc71pFY815XyTnqJOs7nz
tdlTMgDvIKPW0rgC7qZpKlGiox+GTNffzCc+AFA/bD4GW5bp95C2H53ClrTwXhi16cjr3fvE92dn
3UKx+oxDAC6/yYC5nLQT3uDeLKWgz3A6kwI7lOXkDqeQMxOEsCcQsuFA7xd8lKo/WMTMvUgbU7cE
okvl0MsL6VIlE6mBEe/DnYCJfk0zWxBZ4xjMiPZEYM8gNJ2rxjD1anV5FOltAqM16eRm4Xlk1wJp
utzIbL3cKOpiWOcnHkci98p9sYC8SiqofQBFI/WtYa/krJZt4lbUTN0eZkTDqkeHeNIc2RMLxEbV
f2rohhFqqLIVF07SNB6q54H4PA8Mqo+1EPEO+Y80sp5GDR2kuz9KKc237758qroTgXBRcIi/nSiy
3bbrRzPS2zmoKIQVq5YARZjC9g0h4vqTJ2cSNw2uh2EeqPCcmDDppjDTG21xRI2Xa8nQo7LfwaBq
lTbcygaiA58MngW7iPvJdvLAgUzx6r9N5empCyqr61swPAtni7eRwEfx980VZQCjcSVxbgPp1Ifm
wzgdCM14mzQh4dbFUzEn2EGQQa7LmwSA6mcQTnjCQRwFH1dScZngmM3xtdCTxDcN6Vr6dqjg5JjA
H2odragkCM9Xqj2S/1kAwbaMYqO4FLm1kZX+U8zERcTXvNGQZm4OwiRyAvJ1AWgxQ4r8kLT2hmzD
3mzcnlSrshyo6Txkv3wQf+BOUfHozW2gv12RULRiNOrQ051prA1+tfmSqRpjZVHVeDD8myrjfQoI
hbQ2FAOrnoeQTqit+MxV815UHIdjkIef3aWys/uah7Vn+BOCJ/2Vc+TdLbmISRqLU3qjTUJkk0rQ
hmkA7iV6qccDjdthCTUOou77xnrkSlhSJcyFJs2t2+Nc2Xqtr6y2BxjEzNY3quwsnBsSclRIsdAY
TDQ14fm0b7E4y5px30SdfJFYesExvhBj75+ZaI65WJ92H3n6RoFXWCxpNs8VawUv0fQUTJRVNijL
czrpBcnRUvaKHARG2O9szQpg9aH0dUwGR/pehZr5pKlXG6FIs2XVzYjCalnqAxD8R6Xmj/GLH4Ma
yBPaXDZ520gt3SxdTTXZ/29OAcKYbndeomMjR93vBrPvFRlTS6iCSluizZWwB/ba3WIu9Up7882u
PUZFm9MphzKrPH9xb3FdupW7068vx/r36znz4Qyw1oLJ2Opz8+dG3XCU9ByhG95Hie+7lYPdVwx1
WuaCxt9IwkiLAFpC/zQc4MDqCzBAtMgh4at2WElRcnD5QwgC4NW0hyqLvbSjkNPZFU9rIW5uYTum
x6SaCpExWzHOMpFzpBdI5HtprCMZF24JDygNy2nTMNh6TI2Ob1si2gQR/kPBuwy4wWOC84+l3gtf
1AkexwILLVxW+1KUNbBi01yo+feh1KYY9C+798Pqjnus6z7ThZBc7B7GMv6pyIZSRzAadm2pVyOn
1XL7ln4tGjMIPg6XQA8CQFZh8UQasNdpCWyop0m/lOn7v6n74kKgnRMXGSqi2rCkj3q6l4y7K6wy
6r5kPe9ZpMN5XdBiazUuu0vgAr/hsWDkf494966unb40mfdS/yxqbnytqU0LqfifGI0Sf18ljgCg
A3xCOq3X4dajYsl4vdgZDrnrZUJm6KBQQb2PNTHtFpihR1iINqbiEanzn/BkDnmxqobUOxlJjHuM
ZrOz2Y1uJKnZj/UD9GtEPsYmXqxzoucLwcGvI1znG2yAdEm6eRxe26iKq6mxRMD0Ltqxaa70BCf5
z/Nd+cY9/aWJukbSK3F5lRGXip5Bk2ZfGmszPH+f4g3Fkzx9641davbPoFH9FD/13aRyC40I9aOg
/7jLusreIfmF0E/69EEIbT41ue4oFe6+RnUGRnJjl8VbHlTA8ZJEZ5YF+wNALl8nLpfw8COtlgtp
aK3EpP+W9+570cHn/XkEPCpLGQ9rPs860bNVHhSIpA2sF7Q00W8xtPeItJbJVKx/B/mtQNDrKQ2C
mu93c+nHymkX3S95AlmTKQjQdd1jJcQCw0bzyz1JPzRWrvzQigtzQLhORVizNXEaXXAyPXi3EPN6
8LzyG6dS/cPYOUq4ZiXZHqxbT18e+wu6trt163n4OZqPWRCv3Q5t64gvi8rSWEFr6QKYpVyMD0vZ
IOONllWlUQwvMbhdE3Y5bLEK1cTtEqXTwXuCY5fqNDeYYOSBBa3XNZPZ0DlgT0o8FnlB8ti6h7Z7
gKzAiXs8x2iPtumSfDU/a3eCNL3zf+kTz8sjxftj4m/G+wS66CxRcG1umCe14yMf994lz9yl2IJd
quFmtAfEB5f7h3HHJpB57P1lFxILIwuF9VxMDIo2+2xO5d3kqD52kISQDrRUDDC1NhyWN0AMFG3T
8PRyypZCG2PE6y2sHABYAFGlkXhvhqvl8J7wqI+5kijNIeE+6ipOJSU+kExF8gy3J6GlJY6huFL+
Ue20KqeC+SN4YDNV5xUzKaqI+hoETTIJqTgAQGulzegNZi/F6B2xQl0v5NNmzBX+3FJ8W/VVfkIj
wTD9AJC1Opsgtd5TZ3JVH4V4JBOyjXgs3vaiDVzPsjGbvvP9yCerV66bo6quuNBkdYBP/zMYm9Ul
z09hFU4OBT3g+PQJ2RfkG2wadJyVzy9iwWrop64bJ6KyJGWbx58u/Sgi0j3mi3md0vuUoFRREXL8
O2PI/VdGgfdNt3acKhqKIdADix+BDrxiFHlg8sbW8OMS/6TMiVg/e8qNtDb2LR9OAMnk7xJGdR1s
B3YxABGEblzO3uqgICGUHBldW+Z6h6CqSFXUMS+hf/Qzmb7rSPjbwff0Q/jiT0V+6Df1oYu+gmed
jyJ9qfwbHR4M34X6fXZmseYD6Lv8Zl0iT7WOs5COG7JtChRQuK3lBAuZ6xrW982fJXhjnuC26DcE
SBrGsZu9l19qZNYRUYvhN8q8P+fiJLPVYnqC3tdOOp9I8ZSLCB/mOq9K4p90cfWWpZDozvaTtBi+
BNe9rFAJBmQ6jiEBJbodUo5kAQp6TTW25la0LHFh/YpvP7mzx+SiM4RV5aV9+fLt/EMJA5KSKFEh
7d1CeiDCqO1dI7zIJkWQcVB8PRpP9di4utb4cxPTxe+VXA7oSMRQ1Xh4lMT9zhEbSLyxycBjtEMv
SMSL2txjxBAdNvW1WDSDX43+ZwoExgTVmI4ZN1f8AuxKzkWV/1UJRNMtz4typG6ZkwmQr+q9KfpB
gSw9c/NNQd1Mbz6hZ1joQCiWGMcoD+hZEpakJanH8UdGd50e87FnpdKSYZ8FJYDfm5ftYcTLQDoU
5FFDneOYBfTv7PIxIpVq/3CZ2YhVVq6aRyDjPm0e3ltaMmHZEUNoDciMHscWcv3pLQaRr6f8t/wN
arhOg7mJhpqsdTRSM94BwdcDUcUkn73UzWG0x31DB55evDBnJOX9Au4T2cAZwn4f3uP0tdV50CDZ
fvoSb9M5NIFHRyNm3xSXwYnWyuSpKpIcF/qUothUGmF4pz6VhIhva8v+4YZQCANsRpVncVJKP8BK
B9UbtEADxMgXbxoPd72xYDmC4mAlRwH3enJPGTztdD5vcI6hNupfSqt0cOBLjyu21xCpDaO8i/ml
qIiKFvPzJUwHQoc4UlvWReTg/Dazc4uQ+r6Pbd1OSUyvM6PHqIoCfinQgAYbp6JM/WV6PCBvrF80
c96igJYLKagIKen8FpEkY3HO1J/CZqhWr0roJV/TImQwuaSIQOfmbg7tJakRLvg11F9JFRgKUMHf
AQuOnATuWpen3w0qwZ2ltSEysEIAU/CyHRMXGsf8v+alUCN47QgiaAQyTMI2QTjhab0GG2BleFQZ
KSI0yoeDrNVbX43EKWCJ2TduSdY0b40bhfnF8DkxZUjCAYVxNUn6tgrfV7Y8PH0/FUSfyL3sJOCh
2A6XqbgTDAk7AZ32ehmY+HfL9epCvaKP40hqnfEVkDH8BqSygHtzVLZ6KB7dSpI+mtZSo7/WYRXB
PBG3E+kNjTnpA6xryVQKY4N08eFjPKIDt/WePY1qktJQLE1m0ALKYajdFkyIC2eWTYdmQbWkbjYG
hLa4kmGa3fjEMd4oujXH3j2WPrP6rUCgx9gfq3NBUN68isySZkV2Y3HGAedycsawCFtUfrgnVPvH
2fz/+GPHf/5L+96pRbC9m+lRlWA2q0+Ou6/84id4jg7o/bafgTpHdjea5XL8T7eLW1AxlmHmobiY
Av0YZkCU25/y0ukcGmUYKRJK3cO+DjDvHyoJCQQj0kQEyj/jZaFd1X79gVvPfpHy2Oo+gU/Gg78S
Noa8XTiWteqyo/vkvsIVGiWBwPppennO4Yk7k/xWZewV01ghDJFgceQGSPLpIPFAdyUJ9j7CtUwn
Dio/eXNcl7plxskKu/SPHISlal/p0wYiZBU34QJi/kTIozDuIEoS6iv1EN6sv/90RE+jm+OmV7vA
1moeQvhgpRld0A8i2eE+ctLC69FN+eWTfNvyiJQ5xOYRjSpkR+KtnofRTCZxBoufZtpyTbbuPU9b
3ptbwxFtr1kV8JpbI+wzSbmIhKKICaSPzmKIIt4S90z538Chp0mJM8nHt8grsCLSUHlLGSjiT8lG
opUw89PSJHAyAid0ANEoI75KCIhM/GLMFJPwJ8SP/7HXofuXS6ITX0dx16ekaVQxNZsJqK+gf2I0
p/zui1TlkqxMLDNe5ejbcczKaLIUq8szydXPhy0cMaJpgTy8FaXARQUhmK0347JdJHRMaOaezdGw
Iebyg4psytcbk88sfAvhqULKav2hark4p+Blh5UWkWaTXs/bkg4bMybfTSca8F/bVDolcs93vhHH
zwUO7mBC+EvuhFgybBaSvaQPR2/jBuK5lwifNVgq/uqlY8GSs0hmccw5+3wFcu6YC5Wg/P1MCWyt
v9CoMgznewFt3ghcD9tN/PEqyz9a5Th7OAxadAxaot3Kg/8w9/SbZOQLf/DqT1BuPft6jYlcfpEf
uLLRP12+Dt7hVEUhbIRC/pk7oJHYcXZn77TPk2Ur3BR0h1nwEw7TPEAi/o381qeG0PXZi4XXalk+
2+dUoVP0HBntYQr9TbVpKjDzFa2Yhj9trK/QIAyfKF7sATJJLuwIrdr4hk5BSGSk2Z8qTTMURGdX
9GG7OtoYj+GRPkOs6fncsCAClbpVp20EYrXKf6JtQXXzCTpF76IQF5berUK8thUF22166XmtIBzg
NxL4VMZ39i6miH/V56DsbuiTk7rcwN9b5P6cFxuhxMvyiuqmF+zkFFW9PflooCL6G4STMZ8yuTKY
MhgNJFRQFQBGUMDJoWqbsfvLSWId3WsibaXlyAUkITocSUvag1bbn8fQRE/mel7N3TQdGI2tecVm
Yim7LabW88HDJh+6iXrIs0N87u5bWvS/24PTpIMFnCJM1Rx4b+i6kdnvtFGETfjOGJtJJIrj9EH2
k4anWFmcvNbCFjh4HtP3LCbEDoa5aDDv3Dk/Bcf42mf0xmjGEBYy4khfokUwJAlZ/dsvDqYdmX/d
Yc7L4hnKEbR3DEd6vlswZi+xqZ5CQ8kTQuVCEFNEYeSUUbVALJ9qiyIywg2TBuN1Q0c8l9cpeMuF
0LuX/fbj5z4GoCDnqi6Q/VO+fLknmX/JkgYAUxEKm6xl3ID7Cjbtpi+nqrckq7ord0nOO/04tVmN
WZDfs4j6b5dhlhT80lcTU+CVqGqP9H01/q9wgJtc+Bhj2RMpQa6LjbGOlyov855zBVHLWby8i1tC
KPSsTXm/W2+b+sks88IVUQ2Shss7ygThk5ANIYxMwNHrOP8pktvOJMAIZorIARsMi8SXTuqzBFoH
cO47KcILs5TEej1pPOjprDKcJl93ne7Uh03W3/fvYJKgdY9Cm8Bq1DzpfrzsW4Q5jf6bEDzOMuIp
ItBUoEHg1nQp1GeHSNV+KwIonGsMKSXAwalygiLEZeQUh0Nnytl8Kl3p4KFVtSCHAqAMoowfUeBN
3hus8Ww5OvlfX40rb9JoGaTAunn1T1Aa0K9LudhKpGaYbkfV90IxbvFPuMtSrtJfkv+M4HZaRol5
aGYaCUV7vY8uJCrTHq66l4kFc/gocvLDZLusN+bHvphwWrXy0iernULHzsAsd09dbDsZKSOoy7ZX
8F6Bfq2a1wLhR4HRD5pAYbfGUOvgiKwogA46YVo1XHCw5MGCRyLskko9KZM1TwYx7FgorXruirz5
SJUoX4LxpyW7LWUtCkTFFnYmJLYcya7aOhrPzkP7d3Q1Ki9BVpoKoobImAeodDKwQBWT4o6+pz71
/Xg3uklur0Iz53rBm63UxzC7I0+fTxgm83VNLqkP+v/LeLPUyvoYTr3xhofNtlSkWvkPrehcpPzf
tcv5bwSCpBCtN0wRQubjOslA5NUWMfReqtvn2ZNAG9wGwyrZvJ7dDkVNdivN+BPuB+Y0v256s65t
1rOHoRW8/LIR+LJEQOxwWJREsddF/90CIX6jjnSDvB9/pvTFf6FqsHtJ6KLhn6ICCRJS/kKPE1aE
oB8sPw9uqkel1BcSELNSpfXhRmq1TcnB8OvVsEGBm8iqeu2EMnWiL3BKutLtaNYqWzlTo/bqKVA7
Ha3/Z78WFT371m23Ac1cL6KAhoP7j6TmlQ/OQhWGawvYgDOrnWVudwTaUHAhOTOwQZzX9bxxC3uV
U5ikwgf+AvnqZpuB32gqd88+p/iqEFCrIIBCJjEdAOaivDKDR/6jS0LYHpR58ZQ/k/3kpxcHuxzd
8NjEPxeG8/kew8wQBE5OZV180K+oTrvzJFUlmHcpELWCBMApxyMnLuX7qPegmCKrhIbkwtUdpvi7
Nu8kDO+7ajjketyXevAmWUNbQONUtggaWhAeHvSFPNRSIOuP+d1Eht7MmBwBAQKn/N2gDjDT6dS8
mVVT46f3sSRRS7IdAKfmyhsJLI/6JB2IbKNvA0Oe+u4pRy6Vb1AF/KhexocUvnpoQWIk/tNiC6sZ
5YuXe/yNOx6arbk3H6Z5SybRWEXonjzKz0SeUcUK6hFKJ2Bg+VjfhZwu2djTVOM3Cyqx1FIKd9qz
QtNCJ8h7h60lhN3TFPG/O6+mu8xrOLS67IY5H9yAquG8bH1CM/2CYIJp6hgO4CTYvOhUm7axn9Tc
HM4vaOBRPU+BAgYirtzxXizgnLR0uM7dVS4l67atB8CxxLsMf0njwexEs7CenJ5kViWODG8CwZvg
CN+M+OIl/fPAK/y49yFI7psRPyhSVgd0ypJAgTAsAFBP7B4enNH5lInGzblMxkEiMD5h7OBQ69rG
A3W8nH5/n8c8kU19/HqvC1LWrbpx3aJBmM+yUxgozYLCX59dy6VGj5lumNe5bNcnOOwOSQXjNNdJ
Cz1aBQm7eXaaOBT2LMu1ZlbpsgwRwYvmZScDu/ThK7sGZuoSQckIYjd9tzXswv+oSXZIu321fAMy
moNoGM/hjOgLwz9YGpCdgoJOd2svOLSC9ROXnuDouR6CiePDwcV1j2Sqx/n6fwIfVxEYApIo+OXG
QTgYl2noPeAbMzVYK9TBSlmnQsaeaLG167rM1TJLVw3HWv2u7UeJ4e+z5Hn80hJYaR4Qcfczyvwe
DkyDLjC3XDOn4Erxno4zjaAth546uiMKXSXln7/2bnqKG/PUDcLR9b8MO+HvhJAchhgtyWCDNzE5
au37tAacz6BbkpR/brMeQNrwTIOAudihc9YXppyfgVpHYVvkcafmWGJYEPEKUcHmeLWCNWHgCI+B
Irs+kA+ieUXq7HMoxfdsnT0ZtGM/YUzchO+Ket//f36WbzUYSgUSRkHKFOoKX9mQ2aKJm7dhPGfi
vjtAxKEeROx+w2ggm2hPX3BM0kZHESp/+zD+WUk5ye7mkms7dm+9xcdW2oJ5CaZthp2O/GXYsfS2
g74/9Jrm58Y8eTuZDOKhClOQMeq1uZabWQzE95othraNMYY7s3FMPFCOjUZeOq1mmT3YicC1Dp8a
rqC3IgZX/fDBHchkV3tk7tIqKgtdYF4kmHJol3i27j11Nq7CWvOLay5q7aN/wHnm4ZjlCypXc865
jqdMGotn6pYd9vGb+VR8lSo5Ch/PYHGFadJOq6JOpRCGY/de5eMx3OvsqZb9ZeUCu2JAVmyv8Fby
fxuuzWZsJrBqersdLNeDZa1g1wWnJnNkRBgnOkdEdiSHE6zqPsUaa0NLidVoRwkDt75dm9bAXa0u
zbr7Wy0slEpFZFydCOB+6q/UdheHjWwqcRpx65TqP38W/XoXsRRaqhbNS1UXwa2CXD5V9vA/SrdP
52yKANI60ffErpTAlyQdIIrH1TAuTCCdGuB2CYdQVEZxhJS9GocXnawc9sfxiCEocQulHd5HjwXn
VN5Ew8GjZyaSM5ncyjTGNDWZgJSFsJErzSHGgmKot/ypo3w5+NLrxwpSXY10c0NSpSCRdofd0Ars
bhMuktB4Bowkv5kxBMV1nXiSPL6Pv1+AytgHNshEbvQx3Eo9nc/uij2po6FgDGfE5FO+UOnnjTUi
DzRvCK7CH6uW9cUneO5k5oqnlXAslmvLZokBDoSoyi4UCHVcKiwcZYLnCOiRS4pIEb1W1iR9u98z
dVBlLMpeKmXwEMI8JCevOsWxDPstCWav/HUg4E4YRyd+3ZDz06O+l54kdqZQEIYdoTbBM+nj/2fR
5WOXD6uc6E4s3PSqvgl04y612p83giRVGEBiT3jPcrzPR2d1ULZorXP2oZaHMghBpcxdnrbJy9Yp
BJ+qzkyxo+UFrZKez5SSYNhNwSAOIGT3vIVBIjadvkjPJbKb1ksCYZJTcBqbwPW1olzRHkMydLSO
ncgAg1VsxIMh9sUVXoimAtg4CY3qdBU9S4mAQEOBKrMdYP5gpMYoBR3MSBCbl8RuXv73HC8XdsVI
o7xzM2UcbM7YG76mVC/piYqoul1e6Qfq8xZAjL2M9yEeAh48q6YOkQDjx0CkHTv/9S90iINlzjdn
+I1tAn4ejidGuW5wyVwFTIfozyocAhAy89b3gflxTPS5M/EXhRfpwp84MjbkSPtotnNCsoav7Eti
lFQHnezhMOaO2LvR5AdJQYJ5tf2r2tNDaZbQ2nljqeTk4VK3TCQflU86zfgvo2BsWDtRtF9JizjB
CqeGLOmYXimZH47ClOxGIO4RHfQl+tQWltmsjsjXbWR5dGgRlQRSbTvRo9q63c1UxrkTvSlyPOKW
sf9PnN9QI3d8M3arAdQjgnSndOX3h1wWOzMD6Dy78XknkueuLZsXi3dTElcPv4WlkaG1FXnbP1vN
67y3an9BWUu1HAhjdvVOxSQuK737X2SGkMR0zv+qjENVxSH4I3tCHyAOdDcdEDDu/RIuy5ToN6s8
rdO1HI5JJuC/XZCZjdmbYgSaYVWIY6GL1zlw0gjQdZ438AvD1hRe8x5Siy8VcYVCavONMJ1cN6zF
puOEB21NY8+YeJNxaMcCL1OIsTDL/P1fZOXcbCH7Ygmxfupp8hI2MbT2gdwQ6RQplsTYGl0n1REW
72kPWdysB5ePZmdt0FPb0QzRqWvU2w43rJ82AUOvMj+TnAdIQ1ZVZmk9RP30P/ePjtcu/ll/cXK/
N7Z48m+d8jhDHtn1faTtabHGhtkzhdZy/iKwWNUKfoIKB3wk8gUDDQoz1IKQDKI5W6N2vcobAvUc
eTE25o41kY+80RgciopL2Ip9Oa7DDRYHdB4sZBPw25xVPX7RScWL91RI4ugpc5QN0Ja1jqOaXWzV
2IHg+uriQR9bv3roRmU4a3Rq69ZPpdlfx1vakT2sTMomlu6/Q5Cf4BpzSBEE9n6ESjmxZ0ft0ymR
IFyLln0THLE1uznXRXwAlvvzt0tNY9uncnl83XKFj9/SVF13fgw7+J9yXNiULCQI+1hyMHvUNHuf
rPg+G7jE5xcwM/2iLyVhuvBFHOwbQseekQ3Oxf0q+bv/R8uCSFkhVRWB1u4Ub29ILiEM14h6tHNn
VNKZjcWhvXg5Hi/zw6PGa34lY4bdiQrHvNVb+IJU4aXlyloXAt4dEqtWIT9CKvp2102GxC2hVTy/
frFqbcrgu+8G1LihtwFWSZ6cZXdhVWQ4MTfKmQUMBd0Poqud1TIRYqtpiJwHyKU0MFi8Lq9/Kc7j
Qdo0n7wB1JJQdI2JkeLfBQkdsv1Y2Kw5MvUBsLzao0sq5GlP/DU1hsVJObZ8fTh/IgRqpe/pbw43
VQgL2kUESDjReant2Ll9o+B1Gb2XO6DhiazjEZERnPbr1oSHXsIu6JLUHngaHWn2aGdzmHjvPmLD
DngXrPw7P6MtghHOJVvL2LImqfwMPyg4VhY/G6uaKbh20+S8QU1vqHd7m2+Pw592OyOTk8/Golh3
V4rOitbaeVfaZc7Zf84IIRyQA2gKuamQuGkk1vgr/2pWHsKRul/4yF8Lr96NLzJNlaTrf/OBAGEW
Z8/N3Mv1q88NLemsWKtvxplCy/cYMmgHUraMWGEnvuh60T69MzbtGouEEGLWBu5WsLNqKjV0ZPeX
5XxRw9GPuaoPwxLuhI/F/ukrPlMbsjRCIcw7wcovfFU5t4UVJD9Gxy0YH9O6CqZ83NibMJxpzP0i
7qyupSJEMWWa61yAe5W/E8QEeERR8KKxuD/AN5QvIB+fZH/tXt11jVgEjG+xvfh9LtezNOmqJXjT
HVGUAXX2VYNgv2jOX92ku8U1PfNPr0iimhFsKqfuEzTa2ze9We6fDswt1cWD2dq3PsNiAWNGcIof
yLmelaFMUQvfGpp2wy6E1VhOyToYnD4f54r2nW9soVe7urfbIr8mX2oJg+APpbFTD27g99vx9pjH
HIgKpdwN41cTCQtG5S7wkzgz6XI/xweMPfsNpgqlMTgqMbPK2bfKtfzrRvrB0h+m/thCIcaOoYFa
1r0TL+qomrE7fERM2F7qosTw6L0l2GSqgnTbjoz3fYHgNbTy5cH3Q+mjnxZi9WfWUqxY4V8kzsnv
qId9Zlbfwem/jO3GnQuLopDIuLn/NtiIKFB5gg13I6cdA9mMZVHHFmsd3OAq9Y1sh29/9ujUtbZo
c9vwfdmtmS3x+H8xzdY/Hbpojhq5aspQphB7vC1SqnppM36DYX5phGkPZ5d1teNwoat6kjEsDoPG
bN1KoxnpXasXPw1vXc1ISU/pJgHgFGMzwj5jjIgo6xGvmYetto4kb6ronFHf7otwLpm34k88ZIuA
tloiZySsWhNMQN9VEj8LtRZaSkj4ApT+Ofr7KVCWqUJFyOJWoPKgirzaKYxWY8Z4KewFd40/Jv6r
KHhAjrkhEjbjo+h/BrBTOlqkSlaj01OofXz7QiRHHoe3k2xDYsNeBKWZA+PB67BBpv13iwbF5NV/
JxfHR4XmC/9A/LazJh08jLv0HM3/bRNejKYruJbTZ7rqe16LmspFtoER7mS9ygYkvJ9tIXPhVa4y
QCxXQ4//5/8xjZ3X7CBcdnFQd3Yto5TEy5QfbaSan53QGA671tCcqpzOMxgdU6ooITA7VzoWeMaI
vA9jzvjQ7I0T+9U519OD7Qb2c9Ilp72qZ2ihoPsVjz2+EZ3Jmv87PPYbyF7IWvm2AhDxLUfXB5bu
iNqugBHK8iJiCfCZbggOl2n4vuIQXQ87zSx+3edZLOxx+qHoppplHcRfKBLeZl0rl+O2QVrY9nd/
9Cn6YIkawW0KqUJxjh5kO6jJHkugkBGSALl8damV2ZxCt1KvA+NWUvoU5I4DFBtMTGbEFxwKF00b
GNxXgnsxwDB1mVut/YCOQvWFh6A1vLgktit5jY1MqyikfAEPG9c9lBA/TDfFzPYFxTGtnTe0X4ZE
2vLU9uDI/4TWIdwjm0WOjaxcrsgSgeuoyd1OCFRpY+pJ6WJheizfV3dKjiW+BnJPGfw+0l3Ejppb
X2rquzMy9NB+GM3lMTeHGxYaEkCgjVWEsqM9mqncPiR17GXTYon7zQuZiEL5ctOXl5KOk5owPCuw
9xV+oEJihMj+MqQwngiH5QOaW0gDTvBLSCw2wxoLt+WpyUkmzAi9qQOCoI/cdePAXCVBxJ4kb0nl
EFJIERcDSjievfVmcSaQT3xozh3a0FSW/ku6WghcXLr2s6Y42NEG2BtqPhcIHKaYZYAY4DiGxqIP
ddb0zdp1Kp6S0ffvfHZqmQUJwDwfVcOJeQmryYGJLxxrwybOnzE70zbajP5wzPfLmcFxjlmHKLP0
ZZa/KjJ8+swKReNFcpsaVPqXwNES8s8sISAas9GTI1kOnVuDoG8Klr1iVf3ucI4PHOYnijLvxDJ+
rh4S5kaNJwRlRuCTfj+KT/JYKrWWLOQXSw4e9Y9zmhhEXzpcSLxvovdKmctmxukDjZHR6CFvvDhR
7hHrMZGPmsBLF3BaHwqBTVTKmeopIS1ju0EejYLB1BWCNeG2XrOR4IOOEqZ5vlhF8oDr8qwYAyrH
vt2uJM+2rnlybgtObdVhbbK6bgHMk5hUgieP+F+XcnYHQrv4ejZQap45MQGIVIDzsdUCEnfvoZWG
iJ+7KC+NA1QsQO7rc5tob6f9ZAe9WBg2fHWrzR+5S0FGdYuMr+9BuWYDRSQR1EHLHefpuk1h9Gyy
6eTn2hoW6jPU9yFseAmZw+K0CfaWtrin+XZCnOLIbDFL9+JtiwxQLxBSjVDVR0Z+IXqPcNMLOErV
i+ym4cql7C8tGDsChCzOSjjFk7m6pCJWHBNzPyX/iryKu93p0IxX4f1PXoRL66RSdKGA/HH6RnqE
hZcTA7DXEO5aN1xm9TzzkIB6OYOIQZN0TG4kgzt4vGVA6prm/DKbyHe4c0SHs/nvqEBshFiAI9FY
yddlVl85K0uFeVH6wFK0ZfhTTXQeFYT1rszFlwdwxt22+Ap3+enoRATTm/E+6fvdIS79kpD6/12e
Ubku6hwUN4UWC9oGOAG3GBb57PzT9OmKHnitQUkvPQ5sESvBDUUYCL8u1jcMToporc82Yk8R6/I5
a9gBX/8/s6B2waW6+NZ2hGIYqTFZCVy6EMtKIdPfElvs9bY+az439H2vowu7wrgsEVMuBbDI99jk
WEYy5kqKfofSmTm9tz/F1DwF85TI33m9+AF9oQAVU3oTuS26oq/8dj1vwfdABp2eJy7rhDV++WNI
Vnt01fSqdCdjtqsiwXaY55YFp9FVZzHjrSdLb34Xp4HDUhiX7qtVWm58kOsz3PEVVDsuOseC3V8H
3qt8/K2XgBNMp5RjGTkoYI80fPuy4mh75YFCQxkpeb51F0N84ACYQRLFNxSvHCcuGRPRsQ/qkjxb
tUq3yQp3tKcyLVNdsLMiZ+DgCVJ2qtO3rw64ZbAMu8fiMBskmuJVUnR/nrMGaPg98VJrjkj/0kAI
qvfeWpjClDRfJ+VTYj0t4WXxR+Sj66Xpj30mprEz+zsy9jLXrMYKmQgdOzuxOpKMxC3l7qabhOSv
etO6lfFl45vaj8XZRYO9x27Q9Q0Xh2thY0GAkDWQMx+/5TB3+L641DEFLknJ23SimSWhSdtiGfMO
FwSA4Q1P1/tP2rpHdtacpTw3NjeTYYglksOqwgTN21Mj78mXQP4R8V8Q8QWa+9LV5DYeU3kdxzZi
cdkdMpnXe4SmDChyfC88ua+YPC1D9bayvfSZ0Tro6X1ahZQQfJ3eWeKbbrTXS7JBbGkYZNw7ZEYs
NnjPGuTm4j2viutnWpRTSVP4HXzpTyn8HAPxKLLxr4QGTTgO9qryb2sZ159tcEk5Rr3iCTMxQ05Z
tyAnXJlkP2o7hTB5nmYCx4+mJcmK3VXzSID1LvnUdV/edqXZwgncWS8M77FwZ7o926M+kABo0Hce
jnIuIwGTUFgYT1f7ycmjcvlzyje1NezJMDoaqArbYM5ibt3oC4ZD01X5PQsOps7DTiODHDZFecUF
0t8OjBBOa0FgFZcArwI+iaJJzqiycV/hIyAArD4MtT4av8hHki7iMgjeAfq4tJjz38MAk6hOBNCk
+m095UweFqhOo8DBBMhuvzAe+SAl5Z9NASrLbKS9ad/GGehrFJwvwi3183nsrdVwqtt6Bevg5mk6
bfhXgDexxLDJXzoBUZIF6cDmWlb3gQ2StYr2MJ+zDGwnq8WRgDs3oJtW1uOIpstcI5fJMrgR2fc8
SmYGlY5sMJjw+NQDZpV78kA82y9Mp7kYp2fk5/wK4CHVUP7HeNKfzL0H9KSX44ryZqARpvBzl6cp
a5Tgr1IWwCoRrE2C3H7iYNHoQBRbTzshKDPxVUC4VLJFdCq2YJn2vkA5uXQRPThvsaPf69tga2Pu
e9huvmOVE+PnhmXU52d/4zpG2Da+p9KTdVHrUNHUV+rxS+d+l6fKkPMf6QeT++csUi+f8t8wL/md
uEsfqR9nP6Tm26XZr4NNzvNpw8wSVAaK5Ux3u1MxPhEYlzRbGvfmB2DuSqfXrhEsTtNPaTbDCjRB
HL7ohCU+n8oxJ0x4d3aYFUtn1YqGT/bz+5sjtWtlF6x+hRZWzIBQPrD6124p4sfp6MeHRMeDu35W
/oJ4Qbz6PiAstZ6ZeDMtuBn2vCT+UpOf00JUf8qlXoLlIznvZS7dOYjV3yrrEKjVNe9tQ2emtwSs
FGy9IJ/dPCwBJnqFVWGieg/Hw37Zz+yXYH++h0Iwjw+MG41Jj25YH1Y+zLrVDIIYx2YFjWET/TlY
xa80td598KxRy7bsDSgO1HSvaIbSHVo9lqdDZ7zHD+IaMpp8kTtTY7m3Y4ekoeF1yKXA5aTpducZ
bwisEfqLk840cjEi2oywU/jnTQnj1SMNu7tjBd6qLptfWHjdkzlGvHl2fiJObEEwXiFupjlTljUR
vVNH0m7eDglfduJ8HWt3DypjeQ7o6gFLJFCef8fq7Tbdor6EtO7IXGfGz7zujXohtL/HmGzZSGT1
MiRfM5qmD1UGPIy/dNVNhBz1jo3DZSBJcy4Z6MrrYprmedabbbzVjAc9cRK3g8G1n5joDP+YjMhR
lkHhVx/qZxqJmfvmTpOGPfXYG6krJj3vH8EfNSdkf0BJk8HxuGckzl6czQM/P3L2OIPbqyg4keXF
SlfAbSZf1xtalKKwLTHPsNtTpcHuJBAcDT9Ml0eb+DbhjFdD4nIRB6pY1V7xNfFiLqouuVLMZNxY
Rd6E3BQsR5RxwJZ27e2NtD+UptwSc7ra22O9kXuZvjHgOfn+zew36vQmYlnkpxboNHtP8zEnA5L+
N37GGl6vzfs85xmjouIutW2AIDIX/Wn9lZOf22YuYzlnR0UIDiwCAYsetQdAj/7GigZDfFkh+ZyO
/AfA/bwAuUu8tM1wUAq2fYfFNJ2mllROFm9xFnSEaXm5EuQHaZdjs9pjwd2oCsVO7u8nlo2NFe1z
5PDqtcHDtoFtUJlfGaNQaBejWTNUtsunckvllkEbTjJLKFkAYt71dYCMGkj+97+7VmBTNkF+TNma
F+gPMr09ytTwixSUTXCysU+1f41dY0nTyTAGAqQK3UEz5lQrAj4tkAfBQVG1bR9KHcdV1nolniEM
8I49kKA3oEphn75QH11QpRfMnyF1E5UshLVVPp5+6Z/wr5/l7deXHzSur+XOHcgs8kHN5KKTCTej
hA4QazPbFOU1WRhNkbYTfGo1jbMYzLNs9tKDhxcP70vgRq3Br2mExvhTDHJn7AYinkTsl731GsLA
LjQY1ESqXDgxmWfZuNsP8/STED/r03iqXY+vxpv9aF6bV3gwgBeNi4kUP9FFzyIZ9xNiXtTwrUEj
HmVrUFsJjqRIv/M+8JrSkzFyKaVNSxsn5QTwuYjGQGzoiCCw9nGjsgfr3MD66I/pkzzn+UbImbQl
3RlbJrUKMeZnBXF12KWKXBBeiV4BA6QNo2JDxQ5C34896JYgZahSsbudKQkqiWc3Ysvn7pAi4lRA
1YAVDdzXGFY8j4ZQcOfLHi9WH2ImJ7MIuBMmqR9Hrr/pKSnob5c0FxDg4WxjjRUT8SD3+dE3ke1+
jd78TMsnr2fWTn0cosWdfGIkvKrIVr0QZYMhSEIqXcdCkH8ttSROPhLRs1ypSmzdEOr1Nz2C+ZRP
DHUJZy42YTws8VuBBPaL4a/qQYPiqjF7K8QtRiQXx2woOdIU/o4pM9Zf2gc/kCpsVE20OdLNV8jb
jAXG3/+ihJDWSpF/OnLHvOuC2TkxBPg62SNsQE/oXqh9iOeSIOCWEy4PxKJaexCaQ+X7QinQG01C
fqrN5fBYPo1hNb5x4o8q2GvaVT473Mtd735TqF/i6pxrm3HWpCQHX0+askNB+WVifHosbQEymSqT
XAiufHoHuBEgFkKdds/34m0isq16vr5sq0rW5dHzOB1BSFYRi9mYS86TFdJtlElGxFjXNT97MlQH
VUPBUHR6rRxnTS4pbZiTBRrC2rpuWtfVAOf6dNajFFknJgGh+TFIzvp9i//FFAjwkeyDmF7V0q5a
aKGoOqKcy5kmnSldO69ZNXj+/TSPSvDN20wK4gGuzeHVDYiSPBokqJ8N4oLxBakKZKkToWOP5FvL
f5HyxIPPmAiOCSUOBLqtQYG9YzU2hvEIt+GGYpa1f7LMWkKTMzy1i8R5Q/QoIp+4SuvBF1IMUhkY
v5YgLla5tR/uUSyo5GnhGw4ewgHAnUJvV72Nhh74/XtuFuo0WhBtEihUAd0bTXuoYDe6u17ZAN7y
Umf5midLT01VV8JBj4kFwyaNUmfDtzRSILcQWULrJRSy9lHMEgIIElVqmg1OPWM92KWllLbeL/Pf
D8Gx48xds9x0n88jWrugeybKgZ0i9MlWvxJi9T3FZe7jOIPT/BicJD9d5nsEEp5WfysFVzqnaFdR
x9Q6Lozo9if5hIsXFsx0JnsiZYy3PIIY17ZDLlpuVQXArs83rEi9m+JkdBbNObPpcaQIBn4rhbET
zZwVF5u6BgLaNWywaF9+aUwxbNzSKcd7Lw8TtleYiGYwXzvf4/YG3eBHhlZoF3Hpulbcw6tPj4K4
+dpvbPD7TyWPk2Uj3bahjbcmnGrG9DCaiGWAxO5Oep0P0Gqutj0+IHO6u44ivLpXKN9uXGj8scLk
X0TYkpRkOJ6ZZ2diLzCmzOSX7NlXGU66BVqECyb0KEKMaEpSTf7IZ7aNBu4pOKkUYxKUC9CsyNXY
19hAO+e4LrELYL6QN/1BGEpn6lTx8af2vYFN4n7gwXqVbzGHHPig68MzxRpdxnH05WuOqhJKdS2b
3ZN/NHl/sf7mo7AlWVDqqyJVtkMPby+y+ouLBUMR1xDqWCT0uETLEwBDhbwMQZM1BYGMZA24MLcH
piH+kxNPeqYZLO9WjPQSpwdvick/dJyGp4Ov2sxKPtGx5V/sggbiabyNqRSK+LDpA6NujIYBV71k
l83SDpmhTrmTIW7/vmSLx8khCxNvFFobDm7a9WuNjukui3r/n7q6TubmtgfblveT3rDKT9THV5GR
jt4j3f4TF/7sde0rcVdO9YmogE7GS1bbv/Ip+D0SJnoYP/lnRfAux2vQtKZpLkCaCicDiCU3yc7a
cszLENGrHrj3WOj9csQc9r9VnSQ7QWuVabL6Gd8kEy/37vQBgPZ0xZA7Tq9eI6hqMqVF5dIYDds3
EMnjP7Zk4iMqmGp/xAhICnvBJDvsQ+p+1HBxiLwYkZ8vjZaOOn/3bZ5lybDkHcPTBCqTxSm1JwgF
fJXpLSYq4glU1hMgb6MGW6W5sIBUssmIdNo8HoT6AxhpQmCOP+tqScqxBCVbKbwzXXGj/f4gL7E0
KNE7PPrl3AvEW6hJBJVkrLg0KSLmcK2+u7uTHnBUChMSC8cpkm0FO2ythKsSlMMn7K4lckdBsSno
6qPQNqu//XDvrBERqzIq8q/OhuFxOkw13LfcJDZUqaHGP+LXUEBmd6eCuooIa3yVdrprhkdIjEkz
RtaMV2Ht/k0oKwXoDZVjIItthBGvWAbiYhW5DevXi58ringoDwmApGuuvLaJDwDJKM0Cvoub05ub
cKzFJTjqwo5pczMhA+4oMqbYo0ZsbAQwpOajkIKvCTL59b61HhH2OF+jx9rF/GeShqoQuAbuUj5S
iprIYWfRG0xWSu2Q/IqNx6gFwi9XwXlhbxn5BqGcxrAN96g11Wl5mfViNg9cnAK+RK/xz8uFc7sE
JD1p1wLtZnjswbmgqQcB1WOhVjd0MIDEbvJcbqN2Gzi7nNG/FQ9TnIKwAnPVusVZI9Qs4BWbbW2w
YVtFMZHhXX8CEqJYsQN1/azumUagBOLCS2ib42rqtVYzhS7oRWz5mp1uWSCIZ8FHGvnk8ee3U9Vz
bTENXfbbnEUXkMh2vLqEsdU3czVCyNOZ1DgbKWytKrNFPvCh3m2KkWPiaZE6yXrqa/a7IQiQYW/D
7P69ifx6ogHA/UQ/XlfNZz11o44Vs7Syg0wadJ/P4Ocyb5i3AB4FS9TSuGAODbJmHxwgT8ODN/t8
hXPcSOuQYrDEINj+W4yJto4qftVGE3ibKX0Sb2Erlz0RbvmQtrlE/wJO1/uXqtpGqMzDORpo9nlA
W8UYi5q3V/qSIyF3B3WHxqwwMW5T8DmsLZFrD1uTcrtjPBz+rV8FJ6rzcxelA7B/+m9nMNudA3en
OHTkxMiT4UEwAGc3tEqBGbtB3RmC9o394/XQZGTmy/uAkueCATPqBUabFQUdLCY/6BHu0vRTWRLn
8qdNyUGa/ELf1dsJYGB6BRwVDAZFeT6/p9WW9XazX6GvQ87C70WVoz6sYvsMxNO1bONOKi2dnU8h
ZaVIJ1F2QtFzhv5GP6okhS0QtqsV9jpqfEHXl7Hp1kKDWA1QobWt1q5CysbDGA4lcHxtuD3/am9+
FXGzKsdfOYA6AuHHykxWMIHHNqJEg5BS+Usx3R9OCjAfKguIYvfkkJVv19GpTRvTYDcGlEnNy6ru
6/dRRnc1uNFQGhBL3CsuBjHd9bKnBkZHkUloPKE9IPE5HcXk4NUuJNj5DlQwHoYEIMhXvHxlWJik
YiUa3nFDfs/rUBc6AL2zl+yJtVp/dVUY7cLZEnJvheZ42HWITShaUBWsJJG72EsJbH/OMgJA9CNt
Hb1SnBk5e6P/p1zhqd2lUB6tU+kHwACYC3XnpyWSezFvTogcmNKD39rrRUMuaIoObiHKuJ4f4yX+
StkmKITdlIfHnD7pl9gF6MHEEqCR46rnfbrQodr6GfOrlkspTwnrW5RJ0CZSIbdVWJz1V+iXhbcU
9bw1BSS53ARR7aSUwzraqfK7umt/fmjaH91xNzAe0VPhRN15WHF36e0CczdoQISadqLDr/rbGMn3
rBvHsID435j1d4y5/ZnlQJwC0KltwpY1Qw4JP9TLWOf5csU7xjL+nuQuwxFc3KYiI/0xbnwB00oI
yxbuyRIl9UmAmdtHdsnp12r4ngUpbAwx6/kiqfvxvsGKCozQthZSqdngFD6LUnYXZWy2SGaJGeXk
GDkmN822BmoZIrtlJ4g0zt8vCpHS/P2CdqCWqyrpozI3e6YMnrQYp6wLXsvAhLtMqFbsy/UNERTI
ZFUXz2DrtOsk9kckVXbj0FndhoqMDLViVuTJOwIMjU4e6Ik77xVtjfOKmexmAhPr8zg3nkAspNFP
PdSacchq+RtohYb+r2n8JrUbqcQa/5I5Vp4u24rAn7ol1r3XdZHVxcUwepVYxGHByl5frQC+RLsz
z/6X449FPI616fIU9K9F0Bm2GRuzuJygPmpEBArfN9V36F0Klx7ZkEX4W1ss0kWT1LbJF5nXSYQq
K9clqlpXOvp2GTWWWCe8SYoTNY1h9xrZiojCHepSrdaNUQoVkJrqs67KDVS6rKqKc4jxK9ssi+lh
Cz9tnGwOTpLPb1jY7uYSIzAQK6+RL4uFbtsDCf0L6HkP5691VPp7ah3/enIKBq96B+9PXifxNkcn
hRNeU5nMWPD4wTLpLkUGZLFSkps4+TZkp6nGsJajImBofwAo7VwXhv4S3yqazmz7vOgpCfzvygfT
vIXk+UbJJifkltNNinWoor5/2d8vuP3x6SxFmHg6xuj4uU6kXUKBrBNwOiTP9kWk98jxOPFL3ugL
DG/5yaJNlwxWL4oM+l00UeWm9dG1EqaR2FuF0u3BZqWiNJco08nnkd/oh/NAJSmxfKzQ9WH+VFGV
lIRMLu1ZVmM0fOGJ2Cj+copAx63KcZDAx7IAIObE1+cd3d1kRAlg4XCzcLxaonpyNDQ6GFlyvXd9
F6SA4YtI4MJmdJBVU6XcMSshRZjTUE+42SwBmb+hNoeGd9miflFRVsjToRvaH0YQ/O5YoduU77FY
36xq8s4ZG7k+1Os8hzwDDWvcNT09/6lz8uVLVXZbeGWwSX4uaCNY95AbDujnZl7SW/2JwtL2FURS
tBo2ggmHUFSP7I5u6vYjpD1kId4EGGiFNsSCZ1NUY9CfuIqRSC5aqtmM4j+u2amXmjqwSf5mJyPB
5k9wzm5XLFCKu9njjiKwYA1oCNg4jcmSySH6Er0MVSFQurY+gJKilsffs9Hn9fNP1CslED7V2Y+6
uT1sYCcFpSpSC/ZzjPc4Bw7KBeS+TTDrBNPiemuyxuK6rXZH+j1LQ4cqOLoq3f9VgiOOAIAmG4di
/Npj6gynjbfAIt0EMhQvub0EyE0qxDTtobCj6KD9YqWqQYYA/BVsL5/xddmodhdC10jHUiReR8Ch
PHLJQOYfrjUafELRdQ334HwA6PvUGgn3xCoppvNd4kPivfgT3c88rG8cLfOIpLpVvjz36hBzaJlg
GXsxWfSHMRXFTG1wtvz2FIqTsh64Md90++pmQxh2LB43StMWX6TOiRuA5+VjdJ4ZT8EsJLS3vpCo
rvYQq3Pr8gluK+RtlChdiwHLGU7T7Dhwd9FWgOShHG2Y5julR3OyR9MbFjKTH3s5u7OS0CCYi4NQ
bqj+MRciH/109z8A0d12A6kEYLUPNmwbfMesXKEDOYuRpKqaLL+UZNRGUMfw7VuCxTeEBfc7v/XV
i3UVcdfnXQfBTa1ee3dAdCXlMuwG+HYF6Fma5ZA0PMmxLwlQdombrPzbBnaYLrj3UtzlH/rwkMJo
ko7ookHe/2cdX0QaFhoN4f7iUx6TbwsN+6ablzX8x6UOX1ixQSGWmu11vHvkZqLby03W7Q/EoSsJ
Q7ik+M9oLQAGRYsXVv7slhhMH/Y11bfHD6/lUxFo5ZwZT88Vy+hZ6rDxn/68/Pma80jqimKY6tv1
8/m36ox06qx9FotzkWyBRLlu9tUYXhmv3q4ZoOaD/8oo1LQKpaON+zhzmmomLYFe3x0Nc3jfs46W
gpbdYajaKOI0d8U1/vnzPnat/jcEIMrPx3i661KJfArnOdQadVwSUdcMvzy75IqloCrgyu0TbJLq
UTLmlWkJnUXPJKiSe/oswvgjctC1uc370d/0ISpdo1Lo0LU3cxO/8lXnwPVihPwxPuxwGciYsTK4
I0pyy/kfLvIXaHQV314Y0wNEXfK59FcmLe3CxYMOSt6O5/Kk1mIky5p6syopXrqZLpuP7DXTyYbm
f/OF30PQfud5qoKAsDRBcWzpizvE5he9P1OI3AjZKEJcQSVC90457eVbDFb0HUFs9gQ3dKufXbsS
R+WWceGX5db40veNkS7S32CCaFT6cIoxNfqr7OAn9ekrMi0unrqVCqsUbGdMbO/fxNnPvCKQxNos
fVShsSIY16zNVurBKUxJdH+bBqFw2uCQjdbzWFSb1dZ90YJjhar5xCMzdTG6pm3DFrEw2rZmZPMj
AhjMcyoTzauZprXg5i5bg5eQC2tVmzXvXkgIwwmDrJNV+I7dO6PxQQFmFE7OmIM/YZk5cUgEcWJ8
OdA6V+c5qYwx1GC+gxxgwkAR8mILwRX0KH6RTG9yr+Kd0o+IFAxoKRLb3CDOMHt1zb41GbV8TBZB
K1MSGwYNGbKDkmR/KnnI0nw87rSnckQW+E62GXMswBpziprbTwib+MAm1/UxPmaStsX6whnbBM/d
yBt9FM5VZBHktDDEusIec7W7LMu2RDoqPih76qSN8shsGau/GdcLS4VYX2YlSnOZDTuORmbRx4uR
w7EO4/YxZazO2PycJAiFhJwg6zv49gpsVHToNCzose6is8avwpC3LMo5Ior060f0nOsckpaovGJw
bG/Z1oiMV4kVL5+sWrKnecYFdPfZHHchnpefVacc/J3EzJHx+ntDB5iNEzJqLQH/mT3XyrYc8hgV
n3G93SHaeWv515EJ1dzgZJaNQSH8x0HmK6Q+hl0mPQPUWnR5UJz3fYpjahCS8yyeGhWJBzAdyJOk
Ix8VWlmQ/sMPh0UIH6jfcaaX/bRIlpQjse16vcZ14Ngj3jLRXfiTEnSnmczSMD/Dxf9UBCds1g+5
XXwKkanD0JiCw/k8Q2TryBLoJTn/FS49joMphMkr7pvGaey31aALaF1eJE6Xi0UTFJMe/8/8SH5E
R8Zf4eQhjv9yeM7fjmiSd9aZ1R3pEAelEmN0sjYtGHtKAxW9q0FQNjXZaiGdIURdGjUI9yfiU8pN
fBRhX3yUMIF1/hUq0oSxCeUOFBVuVxFEjz/oRaCXuMSyMsmlm60uRQjOyYtcOsayAyoTlZ1o0f5I
b82uXjtD3ufKhzKKS+ihcsoWlotxfoJAldTFcCF1OrS2/dTYcyqtIZtPF64coY7O5/hqb0y88dda
4VJL2HceHyxbkoGFw6LJBjADtn8A0qAJRMgQb5hBJ7u0bvegXTGBcZkIUBHDLf0uj5Bko2BBhnwc
/Pf4WrWralUulfS7M3zOKM8L5Si1W+aJT9mkGpdHCB/SlSgmtY0TSZ3D7pq5D9bilQiCjMO+sdoX
X+/O804FcuO29DEaaPM0xVnoC2+PJvEj6FKKP7Ymi+yGeZZol80hf9JC3XkCo8LRtGIWLudVAoYj
KuT4/5MyYPI1Lkr48kr8ZNeCHkJh2eT3nHQ72IQV0Adz6SJySLt9XcUeDR+OmUX0JujTN52Ot02I
uqS8LPs7gh37U0Pq3MpZhVMNtPjSFznR8N12LlPCLLgCu5XVUNwA7HWjB9DNW8zH6x7buQDs7cnO
3WHb9pcsOXrmk1k2I+yjQPd92JOkXjAPGQIIDknoUlYFIttczTH6NLlMUw2GzdvyCJ0+up/SI7Sg
VicOt1lz/AClSBdXaIHkHrCzpgaTcmsS7gRBAl6sgSGpidtkhnxKvcxSBhb4zdhIhYDoxh1Eufml
QQunbHgpqgiyxlfMhD1CeWxVYo9ps/3nl2Ze3CoOjB5yMXr7JaUonLFu7aSz/UWlHU8ugrbJuSPG
V/axPyEZVBmlcGIMK7MxPraBWDU948TmsQq0hSWIaO6y3BeP8uRPik4zDGQIulCQvjTtIDDvTqpT
s3qTusztPgo7dDV5ph7v1v43Oyy179zqAQZXruY9JvZtSb2XR+xLLsVPhKnu7B8LCjSz7ClBvRVx
qtIVWq0RL8RQcUacHrrmcpliNPwnci60TL6QZ8xymPqvL9bgj+a2qhWS8/SfeoKvNeoWAJ8Uhbf+
Egxe4PRUx6dUg0xp9/chykSH6FvkE2uzDWPLAwc5cdP1mz6YrI9b9QaPok30ymFfdoU+8gxR17qs
XJdqCqJbcqdZ2F+7UCag3Deeq94NbyrNB7EbRfuQLyMMxcAskrIh0V+tKQw+az7myaZ71Eji5Eu2
sKvUpWrFqK1V4cUSroaJfErdmd8MJyDgoCB1pla3pDZhPWZVSkXmKQ104rib79aY2a32lz91lcnH
xVLBxhLaZ/M7iGTJeoPwmtbBBCKSfPyfnd5bLtltYeJP7klRAN4XpwGh6y5dIlOcHHIM3OyeUusx
o5Zn7h8RLWOnMzD5rQv82XV+ZnpR4EigPg1sAxXN5PDtu+WuUJ8bHw1zzSyyPXOBX9dUlGWik7XO
v4IYrt8u9buvzy+Q4+c1dCSw0VF8bxF/Cjkno0i1dgd9lt2p5CRdx343N0L/IzWyO0us7EKXQmuu
KyTv4hYWFRZPeIXeapwIyRUyKb6ldxwq9f78405o4aWvB2pN6AaW+gOiL0cjc+GA5rn9e/artwTP
JHRnUOTPSi7mzRTFEf/irxQUpHPodFgPehriNu7uehxUq8lQEl9YNguXS8AbVEU7uciYCh5YkOl9
OJ7yMgzCeKAYzFJ6TKFeczjS7zocJwdCqc+pZxZAJIehKYwaNnyWugM+Hm07Jl4nqjWTVH3qkzfj
6vy6RpdrWeZKkrgvD859pxZfmfSmPuMZN6XulMAzaWZrouptyou07oeCaa2RllrFzydteb25iGA/
xXuXYNscfCm+wuTRngu2ckVVMUOKof1wDIpk3HTlhgiyRzg8bFuK24ptN/O2Ss2LwQDXqT7EnMKe
QxQG+isXZqii4stzpvd/dgEXVqOjcat8d779bb6m8AV9XMMhKBQwYogjnb3qZjIqvUL09pqy2jVY
kAcXbyCHT+7kFfGi4KOBnKA0CzVcemzXnElp0O7TEHivvI0DXvWewX4pzRIexn4A1xyTm2MVM68F
x5FuqS82ZQglBGhHmfZG6d5AzxEuHB5V23Y7OdtBAW7443IHM+fsGWBHY58J0aXLfN0vfNDInWRQ
8OfeMXxF8Mq5bITzHHi1R05SIitQ850hpvMFSjMR/Wz9DNn+LoOPIRSRBCtfptoJp1tU95WgWE5B
9TknPHpsWqo21olnbrJczyJ3VaQfnoTZkjqTloEOdD3YAbku54v3n6Nl80e+ddW8WMtPG8Wh7kZ5
TXzcI4jJf5W11pM17esJapziYxOCebamMRPDEPRl5NcDIPP2wHzISUYyHHni+zUFTAQgms1Q/Q1J
fy/Z0L07zWGJykRPa8gZkKYFq+1HauRmXD6ZnCXgCatdgQzHclxTmQX97sKcyRtvvFnhItZYPQ79
ZpgbbYdk4+6XTZijJIZ9I4oFZ+FOyefHakqKFCEXsoWc/QW6jeudICMj90FRARkyOrm3w+1sZgZm
P2R/xjxgCGrJ9UovESsKRE+2mUQceGeX0tq0aYrBDf4CJnmGx/QCwrsZFw7rXzYp1VjBed2dhbvi
wiTUXra3LMT7fTisRENX0L21A1CABViBRkYQjk6QTF+IVSAFPdeOS53ZbGnXD8qOk9a6BSgtQAF9
WQiu8QL5fWLXMA0IRa8vAHlrKGKWuyWJuARCd0TqLcX+Y+2nhKn30yJLJoNQSPlmL0fJBietQ3sE
8RGDqnTekm6i2emrFfDub1prE86Li65kBiiM5Cgkc3P0yVunIYrRg0jWRZG+VnjmtiD7wuJpkGCC
vHK1z5Cn/tVZG3APbHWwKYfriDb20s8eX2LYwo2THiyib2NFyqkADW1GlRI9V5BT6gfy5/cAIYfp
yTDSOQeo6zDwnnYvJtV/rVvbWqJdv/wRDo/Ur58fmsSw7EK9dRaZFNYgjzOgdzkxebX2FbuJ/SOt
HmpoRRW6MTMG98dwxl8PEu00h6CsSPbnS8x4ifC06hF1wpxg1SUzlAJLcmc2QHAqA6h88vLTGIyb
qRK0uDRbBUU0gwYXqGSKM/nehmApld2o0ZHhuIGwtvCDOuY5hdh9PCHrGNbLn2oje2TlP5WOqHqM
59P6pltOBg7jRp3VacJod06JHh2SM8Ogz73uyLGgV6+0HirBWCxvMNhimd7lxcbWId2UD3s6wQ5d
8Vtxd07xQXvdCAKaWCCrhERPBAGFwgk5XSo51yA4VjR6GGWoQP3Y7srmDVQzUgVSrc7+eJD4ZrGi
g5Q8MMRS2VyRyjq94Zzl8USOJszME5KrI+UqgW5/CwxR0FcgbVzM54aktwwTGX8BgtR9m5ksGSK7
ZrQx9pyjk2eUuAzRFMieRyOOXOl9p8XMnwMWQNdf7hOSXnIRMWmNYro8daUY47x1gJbKxVKw/HS0
g3VRlIgfd7wz2otdCOArxfUxw6BSqmOkMfQs+dZ40201PXpV6ljGqimXITL4O1qTJXX1/rvk3Y/2
o0Wdz/oRthsJxSVCJCG6VierPI8Efx3sqHvr3T71mW2a0tX7gSVhckz1zPgpLkANaaexJBaMYAxu
0FVVWXYGyqJgSNBhabtHWrYakkyK3QBu0TrjHA/TYQ5Fa0Ci4FaFcUhGDnNZi0oFJ3CtnY7HAtZe
9JLPhcYuebNxVAU7av6g4nyKuQ9r7KPd5y2yCiOmN94aeG29E2yztm6IIjfDAjrNhMeRQhk8ZSpA
CcMauR4bYQDHpsdNrl5KzdiySlT7+APpO5aejwoQisAjdzHrnTotNtB3fD7l25JARRmhH3fZ6XVi
eCnQ/Xq32Udt9t2SD1/I8ix9IuLr5A+slCyqyqXCyl1X9O9XkBovvC0HqXn6ETBmpncOdO2RTsoE
yTdDLFa6bJI+ELnL4TP/WeIrfUUuzB968ZW03oowVinBHAsXcYZJCNi7OdnQSeHekXREylIVHHYo
kdGjlyX48qrfQ/zjnZOywb1opmW/+k2Lih/tuap6d3YGP+OEcdLPHXsNh0A9EK+5IIEAdJCLbZ3e
k7U+UXugXrfStXmatVoFc8B85ElHqyNDHhcxjtBKt9AjRKmVH7BpyEhmGD5nkzhp1RJrmXUqHL2l
JUVljTJmLkOOgrnF9Zil2Ro3GA3LgCYOx/Ns1AMtYXyIrwUpdpi9nzsorWGoJQkRprhZBM4hxHz4
aj7Na/YGOjP26RncNFT1VV9hnd79s4qG4qVgKsZ+iYIc+da1mC1wETbxK8FfQb2MYazv6eEtzBU2
Tp7q0NgIP9fCU6g/7swoAB9aJQNdd9EUaUUbbsXWEh5X7gHTOvStALiTWycescxCYCP769vrCuce
OergGg/HxH8P4dQbAUsSyFdDZ+SQlt4dexOrrmZsFtqCn3IFq+KhrGgMBATShZ8b8XiuzC3s2IHE
DwqdwVEXzjkEFTL508KlCvuP2WFQJFLPxuUQC7ZM3/89eXtKa4Tyaz1zwfO3jiXZP8Bl/MEo8vy8
g86uGiKZRrtk5kD6KCPR/lFfwIqxcxY/dxx+7g+hpUJ3FDoqwBMFELI+Q/O7yHKOx3t5COI7JvDa
IlP8rlMHzX5LRRj3RSEBxo8CFIWHsacecGcuqZNi2mIQMZuQrCbAaNzffNt9hpXCzk8dvtFYLpYX
Kl0CtWUr7yTHas4jzhbCDgSB3ocDZrPedzbH79um1irK+4MyG+8Gipa5OIafAzywMnMb2bcsvJpN
04LxAoCJFuKmewx7flptvUDFy2Mi4Dy0DyOegmLLZme64GjeN3GYSTn3Rasn9CO/bpezmLSahg/3
RyOAPyZzTnt12s5a3T24qJhDURNqT58M8ROeOiD9XzHutFLC9yxTvEf0FUuIAF+zMBcVRY3NGdeR
JZt6g/Jb5G3U4nJaW3OqJImZNOld1OGD7g1twuPnngghKZD+l4n82v6smi5dMwGILyVMYjlMVXjY
fNP5SkpXWs9x/MXNd9g+P8uzDv6zoaG5zoCHuRZmdz0cbuk8KuiIXzWB/jUEvV/pgxo1sU6uMx0s
BBSUnns6bXUQKBbJLmdaAVukOJyLjV3BRiE/vKNAr3GYaVdnQ1xslW+amuhNoBoLRIkf0be/3NL5
+rhGehAYRkKr9icYX24tYyjbLIqDboBRSTU6/SZ3qpSY7FascO6QdIr457Rc5elGYOaz8rY/mk7r
ForlVitfNlV9qcNydpxlLWRkAVU+zFUnE7QZiMlfaoObQ1ZkvaJzRgIKFynhMl1YsoQXukJuhlHR
fFv5clgzMtweaJphhKRob7JF1DPgezdmnZQ7j5FZeBtQ07vP6lZMyO15UkBkVbt1b5mgLxQulkp9
5s0+ik5t0PEWkGLDGjMPvXBVcl/E0EvlaqCUDf3M+QBYBV8CSEzbmbPHR9byaCffIGMyACqmCZuh
jwCSf2UTGRveIBbkEN5JHB7clZeREAuP/KuerJWl9VLhuhM+m2kgRHzgjAZMvdbtWdXxWcx0oEI0
hsWynvkdba3g3FKLtK4AiTckmIHgonplroE1O3KDt3Dcpw46ecXdFf8iqhokuspy00ZLe4C/bs4e
URdvpQervDx8CS/iuwtdO88oIlsVqDaWxAgWAASEvgFyLbaCztt0bext01nYkA44n0B4GRc9Cdxm
brbE0+hOlRMKGSj7L6aMm34FEhftsio4MLZeCja8d2jKTCFyFRGCYiRVAZIsgdRtpp0VtkijfxPf
eAdkbp8BjhF5/3QiifJPfWeCpOiqVecrfngASuNG6gNVE0/e1g/cS9D73FQM5GnqNJenZiZ6H8DE
5sqBZvl19q/UNSzhC2gg+KKFhdStcpVIwrMKidwNIGRerr6QRek9iIYGnHhYxZVkRjQM2Gh9pgjY
BkzNPeugSlgDN3AR52DpiJrHo9kxWqRhn3l1ZVrAOQiuqj/LIguGOfRLWyYp3xcM9Y7hTXgwxnRS
ViWRSi37avBUUQe2RXQH8S/p5bYygu017Qo16cAC/HwiwO36bMJV5WOeWcQ6kYK6+rcayOMyzz7J
fTsUeTSe9PC778x3IkJVdgqVM7RInacjIx0hWEiPEQyXn3az8yQaa3yb7U+UPKGr3J5O9dM5rWDg
UIItRliMwOLSzT39G7zAh9j0i2A7jnJtemoD7tBnTFqNq7uxMoIHDgUZJfmyRzEkogYY/sWIIpKY
ZnK2Ll12ve4zU0JF2DLEh2T8TgexpeM8lpBfiWAAbS3vLN+kHFkGvP5kez5avVj4YUkIXJ3LUsq4
0+PiAxI6iDjDZpWTsUKanROuJqHDiP9n8xftxMOQtP9lEkaoQBCkiikxQjOhL/b93tnXVhT8pC9r
ouDnzrXd6+gMuEo+mvZe5NhXNhkJFWIkDWhdojTrtbQNXCOM78VNphJnhsYb7gHko5r7XK7uhQZ4
F9e4deYtBs7eCNTiu5xEHwngYADQzROBce2t18/HjtSBkVnOByQwG7RNHRXHgcLVgDjP8CYJ7Zcd
XeMcHjLv2OIUtxgd90NVD90jiiF0RKGlbLxQCMg8nQFOpqli1LoCr+HlB7NHjj8WQoKV54Sg0pJa
q6fVUS/w6jU8fI1QHnGWOq5YjIXc02NmeihmgMi6XwmzRsrvsXulYXnmc0IrL06EiTawVFMqjzdC
Tu4s129N3STqmCw6pwiQI98XT9XtRrqLjye4kW4soYQAS6Llts2BzX26NYqhOBl29wl8VsDcYDH/
ldh8NqQPXvj8EYYr1oP2RPnWsmWGTagNukYzObvM/2zdHGtrcXYaAuSTp2pUel48UXCbDj53MgMl
XKlJ6Zi22eWnmoi4+yuhu6O2NLuEGfuXN3Vx8YkwZTEa9MulO6LEPGkLtrg5m99n8UzAFf09UZbl
xaOWy+fjaKMox25RRjF53BO2BNg+798CBCMmyMicuMx2gWYdQ3PxL+Gz3bgD2/qyF2D3vLfJyzwk
V8Ehn/LH/l+X8IcG9QZh2xY/2XG7NdmJuwJPWME2WGh/4UNW3NKVDpeUIAfnTICQyqpzXoeFctEo
yXrgDpPzo0+vG+J0p5TYqoOy3MhMbPqyAwAHQi1bR2q3MhrPHttM75z0ffWmCnFrjDFeaSNMp1ku
cYit745RNp960lVR7SkTiwChb7k5P5O3rjLtfVnpmIRl0KsICw8eIoW7pu1P32c4RuSDtzqr/1+V
v2rHQAX2h1bS9gg7oLiAzz+yuf/macpC+eTdu+25UdLg6NbuyQtXoWdi2sum5Pa+nkq10F3+O3/s
5naXPoB0mllQtKmAjVGKnHHZs2rq0EOw+eoxdwlu8jDb22S4CH623asI6iRkLltwVlJ4GBD2b31P
WebJ6PpaBfz+yFT9bpnNgXKbNQ9eiB8Hg/x4rztt3viRI70D9CaiZRk69xYgW8W2+ofnml2GnVy8
ziqLZEIhQqqLF6E0o4dk2P6twROnFctshE2gTFvrjTj0BUAkNm432niMcZ0nXNWXeftzYPARzKGK
xIpdufYm8+Mlcx5qN6nKLY+P4SvUc+8w3tLYhdE5+vsSVR9r7L+BJ/pT7xnnLEN9xj+apL5naKy2
Jr/82I34ok933dhwVYLDmatgsIzq1YeOseTEYJgw4lGDZJbcBjf++zyl6Dxc8vzlGNYNgtCxIAsC
PhCZXHQp+F5RX4b1y9QVLbLtSpXSYDzEhwzA9+LoysMyuuoaSwFGQNZZ0KiEg/fX4e9LiXkfix1Z
twDzJv0M941rMveWFvTzQhXb0eNSE9YqCXePFZyszx5TEUptcRwx9VvJa0IxeGt+bEYcv0Pwf9I6
UO3ClYKYu4o1pZ7ZUNEqaYWl1RasTZt8Z6R8IZyBH2K3Ps67UzpxBtLANYBGrWoPq83ousXVg6AE
55xytGSM3JefRclyRHWGtmZdB5DGnAhN1Vj/2KHFKhwrsYmKfwuLDrMKqUdXIswmWrHwKajYW/be
Y+AbmWNAYUGxVcWUq/0NHXlGBbBvWGMorx3bE3VCgLlsxC1i+pqjhZiKrhwI33kOtMl+csxm9iHD
ZeGkXTIO412FkDNYrSBJJNdaG/EdwHOxKnc3FtD+lUJ2Hv7CA+ZL3V2Mo2DRxU2yns3QaNR4BKJm
st+KgmKRxrqhSKDNss7U9F8rqRYrP5U+2jhhK5UsRzRVE9n+BonziUT3CtozjrRguQvxis/pT6k+
sH4L1ioIIpVF7hceOMPOgeU+qYGQ5pQUnbHSeqMCPaVQ//OMGzi/5j63s3FqctSARX/vGWocuwxD
RMpYPz/1RK6pXXzdDoJX4uJN0aNdD82zXXH12aNLDrEa/fjB+QTDE8IKCUWYPavGnEm0OIDM5Jld
Es16tieaMrgiRha9q3SMKt5Hr/PWPlyfoExMOamNJLHGRrAwwb7+GEW5mELv/0zH9+dItptbSEBE
/OkUky/S9jS2SqeAdgY/5kHomEWZKr22HwI4L4AX35c1FDqiWrFRskjYuxaz5NuuqJVLD9RnLROz
Nq8npQ+IQr2J0Moub/YU8xkD/yJEo9j3C+AcusIMJdoDFzXzvmzJWvGHrohTOBcZxB5XVJ/fHNdV
nNEB7yTMLR+8XYmO6BCfL5WuvKHpiMJNrzbliQot1gp6/WvcTMsdGPTelVsRTataM0hVZ+QGMIOh
6pwd82W0RDgLAzpky/fLvGrWFW6BRHheeLd+xnGCyvBAergcxzOMylk+DPkFkHCgTrT0tWRo+a/d
ELqgjWSbK3h+TTxP+JcmslaA6QRtzGxRISBMg4MY++PKnEYDtnQobLcx3EcqYJhnKZgmyMNQc5xy
QZxSf2SQOw6F7Ab0ktTGuGV1tYQ5tLCahq4eRgl2vVg90HKpikJXe8K9TPxZaftFsUOD0XDNd8Rh
qSSwJhww5T8rvcRWBvVRonQs4ZHh2qIO2lYyCGr7Rl9eGUpSrAqiLHvRgAO8MDUk9i2KqsrwlXwN
FUqOs9G+EKW47FjNSEpJSjrjaDFEzQdF5lLFvzbLnjFjmiAHzuIosO1vW4JusvaCKis0YRYjC+a3
V3+j+jXWEpElhibh1J4LG7M0QGcSXLgS/mvD6lf9XKBUXgckdcDq2V5c9hbsbVm6SDrVrx8dZe1X
qBaWDl7MoOEQx6o+Sfnl9jsv7+LtKrjS3f4WDBcoebgJVemzug4Saz5A9miUI8oe04F6UwgLoA5k
JFO+tOs89zS7ITQDBaGoUidCeFEn4YLxsB7E4Sj69Uq+wEnr04TJ8CZ4l/OJx3dQDHpO1GypVHbY
ni1CcMOgs0Q64AAn5vnp32oXb+gRfMssmch9AnBgUYypKgqbnwMT9xPLVrVVkhPlJhYuSL9DlKtU
UMHeema3CZPuIMgPm1YURFjwJ99J+vJtJ5zQqEaWiA322F/QCWjUYMAlMVUrGp0PEGPM9e0j171/
qpl/BHobbXhYBPekdB2WhiDwkWkU21z+QiOlhh+cZU7DNFB0vEB+0LnckNPtveWkeNPw8Jjbw9rV
CKoEJ/8NEIRo+BcbS8MrJqSWS8Fg+XOVqpZosWDRKR+XUTx3UvgmwY5GuyjPHayXMFga1cl9vnrF
p3788xfYYDTSxk2wKk5AuNWi2p4/vl0b0me06/4M1hAeDEbV9PK9Nm5F9fzBvUJZN0bMRGhN0g73
P6Ntp8pHEOkNhur6pUJxeCCo+ts6ouz6RgmnHimDxYuVyXYfH1bXGEFNnl0b5zabOMLKi38OPXGg
ZH/T4mSDv18uo7g2TdzDCg24F9wiWVuK/roBx3h0Sjm3j5Wp5LobPMVyoz6+mzSLbf4hucsiaAS3
KE5eQLEluBMeYCS7PT80SJPRT5y7l09AviuWZOMGJ6+aZWT7vM2DXSN/2KEqbt9hip+/o+u/2tCy
6MpJR9KqsV8AWZiW0Rpqr1fCdjdQEAMiuDtYoEiBG5uHu1x1wA/sucwB5o6IhO7PqmHl5rMwma0Y
91g9iypUiw9f4RKmcKgeqImXyOwWvalrO+KA9LowwFZtbifX9OXgfFL50qu9h8vCWlvEv5uxtA1v
J4k6HjcqvnCIHSpdFjh/zR+ihi+PxlL9fudDxNPZleiUpRxOVvWH2/UkH8U9SGESRn3g3Ze7Tx0N
iq+TJf36iPY24zw2+Bz2Jh8D/Hjq3xLait0ygudz2U+Ma8mBb0mzZxJ5bHzWgUK0gCIvKuzht5Bn
eoSrSlIs+BbzcPdePiCpbTWuXPYPbJO0aGEkds3JePLQRlxc4z6fbFx/GdEeClHjDuB+I9CTyyan
S/HLXD1Gv5Pr0NSatdQCQdf88zGjCT4GrYwJPAL+TDRI9JxkpQDpwG5TIswogs4bUgJV8t2MNsHw
o8SufcjUB/uuNphrAHglGs4iEnpUVXROu3Wu9wfrgtPpszJHDyhYAskVriN66Q3s9e/D1geAVKX/
9Txq1IV2tdZRsBu4FEjePCvo801djvXY6QIfMfqCbQGWS84V7zPoyJw9fYOnQF5YJedX+yjuVFUH
c2Pr3l+FOOzyfA7YSq5anj66R61/ed48KXyV6h2eFdvWw0n30uWe2HahhrqG4VNlwG49UEyxroDn
wcFPd4ezV6tTG2vQeQuQ2zmyRH7mrFU1FNDqeFuD78vrEoAlIMcbFFsn4rwo0awT5+0ICBGX8u34
Gn9TjWJQSwJjb7fZA1Qk1FBNFS29W8tahXHjNg1OKlfW522+h6+2/NMxP1dnG93hpTYwvhY74rtt
Tw1ULITroA5X3naF+T8rz8v6XfAKkmqgilHDygEtsQGwjYdeqJx08h8m35a8qqoebSmXxmFFuKSg
Q4yTgJcihJr905idjeMdf3gFRTRTLCEXafgB3dwFE2eX9brAFDqJGLNC0Ppvs9bgtTz0b7NQDW/A
0TE6eLdlHJt1rx6ATK+90MATBBzMSLqLNVba33K4lU6ectqjIl4XjTAcmzwRvXnoigUQEuTPixsr
l6Oz33jQlgrXNTB72dnVsJp1l5pXh0TryLxeiBZ6DfI5XZx8mfrmmdSGBFMVcG7DiskzcriVTA7b
O+Pl2UZNOvREi3CNfCl/aAyti9zOhjHlDTlzYJgx4dfl6+V3qtPXdhMo/GDlddkiHqPFCXFzdWp1
w3VEmQo8vRiBCEOlFluKPhH5r1Q+SGr2Kvo9o/mWv5lK+t8onWviJTlb+rkbP8k0DLqdNqAmE8Q9
KzghYXA2g0jD7WS8VWeqBL6tRfCGJAYoAP7PA3nWjYBNZXvtPWDR5hNU6B1gogZGfFG/VkgTNrjr
vqwkJRYAwTBtGdseE3b+e8QdBFRqP1MycjQb6HuhU30+DgZQCuHMSdwlkI1jJQtlAQF8b7GbDuuU
JQh+q1jToIP3XnD72w9KBoZQneasyzSUbFYkLTUNxoBE/31D2kJHBsU65LNPx46DEYCHHmWC3QI3
LiBu8Z9xoIsuLbYraANP/wcQcejb9rlBVXyCmRtvuTN5+gs4b+jjUhf5989BWh4rlf2RwW4F6Rec
xKwgeyFqKdqnJ0FVtLT8wVlZ/WjbmNgKmhgJePAtMyx1ZnkTScRav5GZudlSGIAI3+LkZN0rUfSY
fyVHPNZumcpDMwFbL9tON3hb1Eq73I2LjjV6C+E9JrTnq3W6ZiI3i0RSLtfMzrQT5jBmEmQzUCbA
Fg62CSFg4T+8JoE0m+4tPZ7gERYqlifhP44rwdfJNDOP0Xs9dHpfSQ5/V4sv7mTFr1guD1MAdwiM
Qo6roUJxFBuXem7aOcJXAydsn3pbi4pFb60PcMWo/WMJWaUc3riDD2yL1p0pO4fM92jOjvmSH/3q
at5ccn/AQ/8jT6VVTVwS5U1uVujt/pE0+KrdJs7HcjhbmUBTKjhRY9+ogZSXawPHIiT/uzLMI2V4
YapGcegNuCJCc1pw3c+M9+ihYguj4bEQI31anTSVsOiaP11k3NSGhPnQFJ+1uFhbGoO8i1RwTb8Q
p87rO/TcXFrfiyZAGpKRfOeDzCOLVWqBPTo+AJFH0MWVxvFLRXiFTtHLSls021mvgX2T6vFdIrl4
Ah6k2Pz+cGhluu9X2mlKmK590jepGLN7cBdedUXkv35Qo1kBum0xWxSKCCrXidkJQqgeB1XvbXNa
dSdC/OP02UtuDQLyvZchIivjzrSRKXSP9YiypmZdDpzFvDQyOuiyapbolU2+Bn+xBxnb0vhZY+fI
uq6jjxEeyASTpj5PUL+YrxcR7qSzqYUN264JUCXiGZfL7jVk8HNsbFj0C7/5VB+alx1tVICDtoa5
U4rq9tLSOEnk088UUgasyS59U3Gn/Guip7TxfRh6tEd0hZQ351p93nxKYM+1ctBBgtYj3S3Y1fwD
3XXjpV3EgEdolvl3UJ6A+kxk9zs4cbauIkLJ58KhWdTwtoa+33f8Ix08bsBguXm9iNugoc4M5E81
cQkyiOjEfBEun1N+23LLBy5BxCy7Uy31+yBIU99oz0+f3z+d91PYXbjEfDsaV1K9ZGRTZ0hQyxkD
xJllCH+7jCf0+lC537MA6+y4p4QPxCvyWahRwgqbNGU8kVhEFsisFrkBjJ5MJzCBJ2EMFZs3oLpb
dNzuZ8pnHGayviNz5C5PQZ4ZHTLSiVfiokPJxjnF91TC4TCNmgWHTxlKezTV6B+Fs5B+XmNv7bIn
xZfam5f+SwlvlrDYPYcJR4xT4fxeq+VBF7PZFEB1iSiTXZZsdKiMD9Zn7AvCv9ynMdo/RAnPILHh
N9gp3YsxrGuVvAAKBEPHdFLq8lnKI7DTfPL5JQpi4QtEmTxkrcoItbLrS/zpwb//R9c69+eUeifZ
uG4FTws7YkiKWiUt7jrIFzM3hyu+cpX+ahZn203dfAKnW4u5NUooaSSyAfk5PPqmQak9jBCINan0
ohbu5uFwTsTO81l90RBNPSahicQ6BkCkW0142eAmbDkehBXQRdjckowYbWlXbxSz1Ix0fuA3YG5h
oqb3/7S1HfcbGCUqPX9Hi7EPzFReMrmMlq7RHV/5oiBJu6CIqjlkVFOVdj947BqpQSNdqcbElybe
B4H6VdkMCluYUArDyER5AZSrb9HQpPVnfv+zIfBGsGvjG5IcLvVOm5XWrHnYCu71HaQrqWxCITjT
cHbLzhGjQBFwDPrfKr+BdxQdUKnqcdZB36ox47f0S4VDa6XcKRrNTT7ZoM8ZUotIucWstsLyVMKN
f8kDHKQg+/h4KmB9b/qRJiQQwFvcqh3ev6JUZk+/AHv3mX8SCuLrSw0U/125NLpYQxSTtQw8Nvty
cAESJEwo8d4PpbGaPQwPd1BDtD7XI4VhEwGGFpgtHmvb1K9Sa2wo5hXBClJ2kxWc4/QXCaZj+mKh
xMzdm2frzcjmp7Kb3Ez+F8jffg4aoBb9WYrEt19DuNngLt5xPHuzBoDgfuA+BiiyurAXUK+3gH9r
jc9ZnruBP7n7Y4hqEZuMw5FcvLyZzGczE7lwxXePcEEEnAMWwpxKivWbwv4JY/XtuA9FbCxsHSP4
AQu1DagtuAkf3X5zHYqv5FlThEiII+C4/aIQrcwkZyyyT6KJ+nStTVFCbbq0nWmx8vHEHvcx2gqd
qSt030p572jPkvXMH3YIQm9bsIsoRmess1mSo4ra2awmRLPr3BCHOjSouBIQ0ifBfCiuZZQMlumT
ukis0dUiUyXAVVfHEWCBVq8ylZVl+9LQqLJNlJ81x95dSDbzKQwO8Pnj5UFuUULpgqw/uxj9rgwH
+MIqYyWrHQtIQ9Vuy0CJ5QHfLGrbHMYJXXlou69TFov/PpgYPsc0coifuTRk4biCUbrL4oPJZ8Cu
crt/70pH6XBJbuPmoRIw3DBGnRcyuD3hb+kDQe5oi00ZPF25uyd39ohGtZLjbV8TtpF1ywgJ0azj
UsAYZYs8Y6o5/47OMBXJkZChkB9rOpqMqqcxCwSGZjJ+0//K4gVo3ZAvEWNjltQh/8Tk/JCCzKuF
k3Uj8Wq42MqeybCxdfaBj0cToLOXHGJrwQ5Czy0OiysmjG6iXMoBcJ6eANTj0HxnPGdHEyZZaKT5
1JaZ0f4TvM7oXBGv568er07XLGVnI8ojxIeOP4fuWNZfIwBHIA1NqaOX+k5B5gyvNAvh3cxG/QpW
uHrtF6k/RniDYQpCPf3Ue9jLbR7Z5gi+ZeTNzvfAQS4evQNwxNQrHfNZojA00Rj1ePHQ8H91VHWW
Dr6JBxzYHaZIRLdovbVJysBb1HoLSdQGhXsetphvOATJvjA47RzKAaebnCxpOjlkwX/TDqZ/IVup
tKddf/63iFvMiEgUSsc4yR2zD8jcEVzLif1JrhohXcG/Mf/55U77MuCRXsD6uaEYHvEPCFkDX4a+
6YqlzBT9Sy7+If/Ed33WqBErxvqNB9xhhCkn+OU9dBkT5dzjWXpXaV8UbFF2jIhBMKXDxzgrkz0H
gSUbNfvzNNPNcP8KOZQMjrFgcLeEktC4HhIZrwLuR1NkIwaTSyhR/gVsV09pmlozsdi3BHfmnkNm
yT2ABNieNFG6MPV+QdD4QBfOASqVIn9Q4uLN8r506aDGYUVe8BL983EAPdLccsmWxBkFZ+DK0CDY
EFSW6eYK8uf1SPBI73rZOz9Dqci+fWjLibn7CP69O8e+H6Q07AqBwv3ZtxWALOEF0CIAzj7Cudag
E+pon/kPS26qtlhdIHNgvP9jmI7h9OaKJ3IXE56pKs/xzxNmHB02hCqM1nQj5sIR4P8cnBcPrLZa
rWQEYxFBtHfg7T4RKTAEJjxckuwj4sKF2Wp37mjKLARZ4i0ybgWC8TMTzpgdthR01N3znzyYyX2V
dSI/uGwi+9UMoBmAdUlTDE360UjNlnsLya0MYcOf2euZuYQpFLEAafvWisvu8kPooiolfblbkJ36
AQSBeLcEeBZrCDn27CdgFsgxYTayG9QmavktJgicwFq1G/FaKCxhbRuSaU4TghWhWTCz4XvWjHEw
PLEkmZ87FZRlc45pW7jOMHe6+KjhvMfmLz9rwxlDKHd0cQrlChM9b+77zMQ1WuWeQxsrleOtoQDW
zKXL0MX7vx1sQEpKDB8/mQ8n1EOHX725qbqGynDHutr2FjRWB2Auqp5nvq1Nhh2plYiQq0dAhNH/
I8fXk+LzKtRsu8+DWwpdQW270fhfZ2XSZ824wV06jhdAj/DaDLNuj5TcHAiuAadiE5i6TSf3bZ2B
LGSizMyfcUxSdczvx1eNBb3c3vW3b3AvLMVt13pJV83Bg3u9JcLQRSTWmx33E2WCyGuAb7qVoPr8
Jl/QAVuXrDguPceL25c+lfnZ6AopYUsHIh+8DBWbgCZaJ9f9oBArOyOJND9c9ggXgPZAN+d+JlQo
hM3r7HgIUpzgP9+smY9AZhnxHVN5kYM/nWfPXVSPO4oPtZetV8prPYFlaCju7UdAok28JiLLR02P
ED98DfsYm5vvvhMtyZ7MzhOitpiGLwnwLvL44Jpjr7fVWeF/2L7itZv3mE/Oun18LBuOPr5MK8Yo
HIWEfED8AXn+98eBd17S9dJkF6VhxDgEn/4d4DDoNhs/vkMUyipGLkrAFJ4mrFpHQmuW578rbJdT
DIuZPrxDMC1W5Qq0w9aiBdrkrBMCuZBnrFPQy9CebTJYtvFrNzfT+vv0tBNiVBlCzdNbAR1ZTcG6
IRL/E7pMgEc/964rSVcoKcnu6NBW86Co97o1XZjrSncIaXMXk+caGx0yHQC9o8TabQEnF6V3wUkx
fcGhyP6NrqclNb++RyWbYjyqi6tATxxlR8jREOphQ05lVGo0qPQoPaaB2rBF4FHzyPLqtrojBup1
JBKOQKvddZElOVqTUC9W4e9SwPgZhzSes+Bj2XeXgMFUezmZq3e84SvItUZ3nBglfRNdAZU1/jRU
zI91NPqu51kpIsExmXKFMf1cVBCalbYOCAx7elpYS8SP1EmodE9oqLQOWkKQ5xS/a6/LrWSsUb6b
/3Kqvnd0jIqQ0nrhlZeoNIbo0tadGr+iA4/NZFGI4jbsblo+lklA5gd6qLFIllfq0PBp0DQBCtmG
5XUryRUOY5n/NOnCan1ViaiP9QKJVUGZDBy3Mb8h6UIDRgn6cyP2XEaeQy/6AkVM/5W/qW/ZOb+a
aR1CL3sZy9WVz/diH9IweYWnxJqGA6pr671oOs13Z8gj0m8KKEi3rUm0E8zfzQ1hvemgKQxbnV4g
CtgVP1Yh+lqzSGX8LF6qU37GM4diia6Nb+TQyDElSZJgk6quiwH/dj1lKX5REFAufNgbc6jjdM6h
3mnnoirjBLsOF4pgeYeSu1JUQY4qiD2uKPOwx+6UImqpOrU63MlkyDPm/aUaxyoh9nF4/fDm0OBu
vzfhf9tdqeOoNHNHyRZQjTxuCNjKwHPpIhQuLg73TYx4pwYM4pzJfAgwbmAO4tZ3LUa9C8+0b7vu
UwFMZH/Rxcyj/6pDnGo61FZ89ZeGJf/rBjbNOgKeQ0O8wu/rvPti1QCE/q6ZBVLkrsCGgCiJnnGx
agSRP5PhPNyzoktvi28sJkYFDGgksAo0cHmLbnhFjUBHz8tdNL1/yxbbSg+Oej0FrgGbXOUzvtUP
YFv+/VycNhbfwJ3rlb4P8oHedGFXx98GrUqtx7Pfi+HC5121cljzv2lgUckLZk3puHk812RGA8XK
kEw0wC6ui0FkyAuJaxOFf1UiDz9xPTBLJnPihDWjm8CNkL4NsxDcupcJ1K+S+NQD7WCOS7WPlfuY
aB/uvr531SlwL2D0xOxvN8VJ8lXRKl8b/U9iYl6MmtZnu34Jx9iUqvkiubB8vc+PkvV5NCjx9mBM
k5uZZl2vjIFBXEB2dNQBAvyOUsxoFYxNV8vL+529vrfOqp329eqVNueEzT912E8q6pMhQ4yreG2S
EdCfJ5AhaB82WXDiJAtYNCGh7FL1ZxOPxccqDD7YVzmqnIaz0sovqbq8okcLqtiZvP+npRY8wf8l
2DX8v/PR0o2W42SimhK6BFgA0pY4Dv2TU6bs+64Jnvdxp8KtuCgKexGVAehKw1tyToc1Z3phyp1D
nuQu3c08dcW8n8BUj7BqDdj0ua7G4cAJ8unf/p2UM9ZlQdYXl8iRBCZxWAkGtPliIiiyAFuipcl4
U27zGuTOqzHTjZGHTkypr046qz4Eg4aEUiIjGzNVHzHHKvdrfjHC7fnGCgf11SQNa75OvUfOnQAM
YK8J7VPaK0aOvnca3rRMV7Occ2FDTXtZHVNhjxeGRavhKKSfM3zdEpxA11Kajwpk4f7VwsjeYq6X
Teadcq5mdtgVAFPSVfWmtVmqqXFrYMlcfw1oX8clvpZ2cLQWYPhUNk8cNrJ3U25ysROzRrvIobUp
LX2pTWNVd6tbLkPV6UTV22+tY6upej+1xuoYgwlZZn3kBPQh/fVY4Y8hxc8uQDxwAWAhU02V80BW
iA8kGLt2ywXrXIFHit0fmzOs5bARkC9svA8A4og6SLdYqhw8h8/l/GGKxRoPneyvyfl3TTx7hNzJ
jZJrN9Ou6fVZL5qiibykBWU6G7byqU6l7Jm9DpmYjbpj87lcSmJIsfRJA8CPSZ1NJ0VwCP+K9/yc
UlYuW6xECaloN+Ac31gFoliBcIcQrg9blZpKl5PnrNwrVZDNLpfLssYovFArx49ifmHTaoHC84jr
5mJ9zzOTfhz3+ZFMnm+x2KClS1JK6biX/qNoHpBVL+8NlIMtSRa2T3EmwKtCeEL5OYfGMgobTZjA
+u5lEYkBGnMYndXXBr1ae9eVgAZEnpRq3AbK/MUBIZ7TOcQChKDfP+xu7Qpg65OfgGcQtuOVwza9
XC9zNpzNq4M+0slVMdv9u71SNlCtGCQo7Ubwz9BrB3LLruINYeGolc48tZXMryqR/RErz0bsCEPw
QZywGHzGfmcPYKcGrxiO1rhgeZgi2FExZuWmUlEx6CmSaKepSMJ9h1aUEuK/1asog6qFeWtmlKJ+
+7ipiKc6PTlgBMOJckXuXxHHyDwoKZnKqaLRB2q6ZOQMofgaqL5zAxePTurqWw3LihO4mNodzx64
HMY7DvifxUyCqTUgfGCkwDjnnSxWkMPRtpyNrjGoXJJXygQ4w39gpfCDwP4soPGU0PBrUYIo7Gzt
AxAC43PNeIQ5wdlklTLc8E75vKJEOryavjr+3mW5EHfWpLMVsrw3tgorTpZP3hA12sLK3PrWAkYR
+rEF5wnH8CFs19ft3TjbAONSZL1lIdDio34JPj53nUsCxdB4jnvX2ewBhfgPTIQqxJ5IOgxOfi1L
1e7LFynNcZB5sX/2CI7DYCzIjjkI2sw/ghmG0w3CTK/K0dQmrO+qmTLs74LDaP83de9IoW3B8Hir
bx+QHnNqg4haQ55Z4cjvP1y9shRkx959+pWi/WJKio11ZY1X1Kk9LoxwOMuJQ9jNHr0tENF4jnVY
r/dbC8scHCxv8GXEx2wReh0JmnssupON8Y873EOLWVLvh2EOsos76R+Gul13SbSxWPBS6vU+uVaF
WS27sC9z0aqgCyXU4UMpN+OoiH0OKvW1p2jw+aV3nbdMlOc4STaQ9GlwPyxsdC1Odo/x708x+TUW
Rw/f1Hvex2NugGZCfqka00JEO/ACf/UA8jHITGIl2oByoiY1MQdgoAgN4HqEG4JEheN4x1yqwkkW
dtYFuEGFvnP8udU5ITS5bNFnuXPIcJl0EBWw3XHdYstDqsG4wHJeMp8TDpX793ufxnPhOiKAtw4j
X98VoA6A1LAB10wFaYFn3Nqs5BCe1AnzazRHzKaPBOyIlxuPlPq+A+OXy6JUBrWX1kipoBA5AMdR
WPX04gC/mtpSsvgIMaMnxLmAOeIxoeRWY1Vjk2kYgNu/vO2P4bXi3qb5xUqhEijn7WyizsrhRlkO
WQGVtMJnDhrLNX4gwLZshjZ3oY2zBUnb3KNtOaD7OSC+qqSyyWtHukml607+pCW4Uoeaj/vqyNoZ
Wx/dDXQ4px3+oFPy/tIeUNjC5yX4SWs9Lv3qFgxIH1ZqVpueFRYvUEXCn7laQVIdsEnJYpCyISRm
NRkneiAhStgLzaS0SpMAB0TpXQkge+k7Vto6cQhQ0NTZdz3SyC02fvtgWewCGcG6BSNFNJ9G40Lh
BituTmOWugD9BdIH4XXlD9txl43S9i4Mefsm73eia/NC8bg9rtnMP9UabXY8Gz791x/kVHc1acVS
vHnvBb54la3/2P0/Kb5c0/oOKrpk/hbj1R0eB8TFp6Rd0jaCM2SCasnKVzNniRCKwMhOMotpZ40b
7gGEQPRLog63nfxm0LETsgOR+N10TXeBSIxy7B+n/jiZbYu/9ZmqJk011JIfU57w+TosOAJTRzUd
D+GGZBZ3ocmIh3dDZUgSupKFgzFEUaYZ+RznIIeCeTcYrPEMKCl/YJltp7k55gEH3US3OGFWnxZ/
JmuDpgWoyYIt7G+gbG80HzMImfDS9BIfwc/NqmZmecXULxA1EKcsXyqgoaL5O0wuMjsiWibALxqX
Cma4GhY/vliES5AD82j5hESx283rVhg91jEqUgH/biukYwzlmXQlnNAlA5Zv3AC57vFS7a7xcEzy
E89Q8RK0Xl2XWSgOucoc40qyZSnPiv34N5BAbj2/U/VtoMOyn9kaqBcbdeCNmRexYA0jBH27W0T3
3usreXIQs/0Q+10VO3mHIbY36Rv7CUbW7G2FAGG93oMbYCHkzsQDqtYIAu2c1bDdyLAG8NCs01p2
PWFvsfTmeS48XCXa7OTbekS466O8iJLYuIMgj/VAkZqTwOD7P6pksJ937StON9kjxo8tW9GCzCW8
pN5tJgAfCAO94eoC7GydINuKfTVnNlONyNIcNOMb/HGRH/QB2uErz49OeRfkFCSi67gp6uG1T89J
l+4WC2uIL3wZXd9e4z8xVqu+cgF6pqGu9ZRK5uXRA7wX2hEZZ6a1sRZmrTUFO9mxE/FQ0xNqh4gt
h9cqgANwoKu7UixVbCdGay2QtxLEWGUzKnwnV0cLctQbeRGtMfG4qaQ/lfn3nPJ+thj0y25DslB9
ZNPauQbRLp6RkZSahjbKwdKNMf29owwqvFKUwmgNpzWo2nThGKLTfnbwLcXYp582MZLtR7HmVUFX
4vMLEwh4D52tbCNpMOhOEz5JxaLsaExLs7qbwyVRPdgRBqyVU4cN0Q2hRFIrz/vvHwe/6ui2bPYc
FaUGSL4wDtvC3ZCo74zafXlxG8JZR7sfpFPs+7J+gaMXnj+x2is2Uk9CtlLpee34WTOPHiHHohWt
wY1Yy1dkC1lggHJJSqXR00SaMq+HCb3qH7+TW8yJ0ooA22R7IKOy1/lJCV7ga/AIija61lqHOPKU
1nQcsLutCQZoLGN7qyBYPxKLNFk5M6OLye+OdDiDW0bMgRkquioerVIfbztwaK7gWKLlx4TxX13Z
N1KRGlWa6vMDsy6t4rZIn/uQit0vFLDr6P5cJ6no+BuHQWXdGEAIN1veh5PZybLaJlxg51ahDdCJ
/bSdIF0HTOzgJxT/QPW8TzElA+T0CIeDGIvYX6uIGD7CFQSSEi98/eN6ao5utIUQ1HoeLqO2jnBo
4qA2GqOx3c1sxBBFJz1DZtcsoOSvxsNOuGB6vSekevFlKMGI8TB7PbyjNLV+vYlJ6Gf6l1asuGGz
z1cF56NMpL+6Jj4ryMyWfbm6d76qhi4lR3hZoKPiXoJ9MQp3YHolHqbEgWvpTlb9Ps6bFbfbEJy2
Ov+ZycvJvH/b4QwuZFxrU9udUmuVCNFPbHrHsnv+ax/WW3R+aTjJ67ENrEcc7qJvPJYyeGf2iWXk
VsRNmkoygSzHwR6lun8Yny4ceq1vsXQoAcZQ3fRY3po65NzjeUYSXlhnBeuyH0EnB3z4AvBKOr5q
QCTjIyYPuBpBd7hFv8gZn3CW44NYV9Im0uVLSxMQSaGSSPcB5JaFVCyKl1Z5Z8f7guCp5qwdCXcf
Pvnk4MFKrpRjdSrw/PCC17/vbM+LLMX90w0tO0IVPoKIQogeZQhED6pGDnzhAEYKvPFff7UzCHxy
0kLzL30n1zMqvQ5RrdcWQWpZdDr7HpJXUkz4kvANCQ6YwF1/ArjvWABTvA3FwyMa3EEd62xcwzdy
5YU/TMAiIIyZ4Rsf2VfW3ENgjuKEJCPfQr0oWDm6D6KcEL1nxQPvKRiyRMniPwbUFOtaEogFyBwj
5NqOoRCDSruXHMQRq1YjSdbJ/gUOzpkovfHgbnwqhHXnALjJlHaXtm3sXZCqgEOd9mjyk8JRKYAX
P8fPnr+jDGhsN9+pU8yyzubYZwPc6A8JmsZeaJzZHmEx7NMqAAL+k8ud4gbZTy1Dx+CTk9CvHCNR
0tx5ZfWLRvJQgDiK4Vbw8ugWUEv0FPfjLSznJcfyLo8+9eLPzjm3QOs/3Iyk48UYFquFvo7kRW2S
4QzVCQ9bDHFK25F6k+WUwmOEoEFiv596gcZz81ZxMHWQzGLrhKLpTnmCZ9eUN6W0Af+3WDbBU2PN
RmyOMvT8OpJ2O0HmJStJRpTqChfIycvVPZp86XmRtPWwMtq+ylNwvUNevXW8iccTqvNkfDm3oXUg
n/uTJ6f02jzZqSA0anREQoNwP7fXkS6QJ8gSGYFSefWE9fpdNiC78yBPS7hE2Wf2qTSbjqdjR9UV
gu1Jyn8idkoBtFeOVI704+KoWLi3XCdqvc7gpALlo218W5Y3lyAm1kFarO2E2+EfmvbWCh6T7msE
0drHRdbR3brBpaC6pqA0i4O9xWB7b8lETEOR6rfbR0PZZkeC7InGe/+ISlIPWKiLT5rV0UbKsB/U
fem6aSzFr9hK/EcgHbBMCPqixFvXetykdutGlITPCttgE8l5JI7PSTV5onGQS8Dr2zt3D9jqI3ai
jg39PTbTmsj+XN0EWiCm/S985o+LZyMhFwTbQtg+TNS30bUPx9txHrYenJiCkIb/m0DoPI9dPUVk
7nXHK+xkn3mt5Hk8bx3b9I/ZMw3Li47gvFRhHcxTfoiPt+XfemDZbDuOgWLI5bIxcx3O6W7j6vGb
XVJPkkX7aJCL9exAGJU4NohR/hIWTddjFnXfwHlTur1lcK6xs23fq7B+ekc+N8JTE3lqHPPaKUUJ
D/DS+o+KQY+MDzU0p6ZEM1aU16oGWnSe04bjCk923wd23zjQ9MwVfvZOLUIMomOPn1GqN88rl952
OxdT7thA64bJ3NzE552ijLgMJcR4nCRxcfH7quF9Dpk3D+UDrzKbO7VyUApRIxzLgFvTRSlUUk/R
nRlI+VPX5fScCvn51EIWReFXE8kvyi/eHEFsabkEEoeE4GRCxYpfectSg5Xqw299vSch9dWBXFGL
0Mu/+KDQEqSj2a1GHvC8LOUmPEqB2N6K4rE2qyy/2n7Y7qF+Rf6H2mBVBgaq5pQNHlj6dcij59Et
MZk8jQwbXNgHgUsg5Jz1ZYQZQZsCPlnaXWm48OMPeFIh7h8uLCdNwepYeHHf5v49woS0lu+kxeB4
3tW/yQrn0X4fHijEbxn83iB0MFD9Q04NdbPNvdwHn4XTX/2NIB0x+KPYfNFGkN0QAvlktGnLXDl+
8x+JPmB1koF5i9j+l+WsXtXPYS0clq60iGaIG5u9I2BetCyUlfwc4u2oERSrNazlQV4+FpCBaWhM
WDKs0SrTLIAvMGrgLTYkSdTV4ENpyL1dr/S5BgmbanDlG6A3epYD9ygC0dLoj5d6aeJ72WeJYINT
AHzPlewp3rF1CbLht5Rgz3t5MXvl3Yx3VAEkjuUf++u6LcWflVHl+4VplZNCTo1bpb4MDeprEPIU
cKYeOdd9j0SgkVToRe3BwXv2j1QH2JWaTYYWvgA0nXXliw93sCt5adWq2iHcfi3dn4pzdzUu46g/
yA35FwIFOH1Z5RRtiPDrKvPkvzXxrBcXVmxIfhYPcRt5427uX5JlnFVIU6yulcuAvhj5agwKS2xA
w0hF4JkXxiAm0aYMmE2D9Rgp6SFoJ8TaYPiuGm1RYOppDmzIFNxW104Ht/rps8T1MDH4LbDJnZ/5
3mwv4ALpFSp6piYmMIKtzB0sjBU0peAEskztY30M8ujXuxYRNRjeJGIXBtpQasywPSBEXek1zThG
xd2n5xPg5TqXibnVc5MiicWO7qqiDoKG7+D/x+gHNgyGsS74mNKlB/7VFhnZltDI/f4i7UqKKTa4
zt0hKQPGFBoUJXBuZ2VOy2652H61ykkI9Z07VtEZe0uv9n6FpRTi2PphRZu50n35nNsrr7t53YOE
wkKPOHG1LI8qebR8NnCNxgOQeRNIW2AY2X8ovTg/3rGawinMBdLfE7rJ75l4Z5xajkvWjteQc6b5
daezbg+XYmdm/4UhCkmf7js9H1hKyP9FA4AWfEvibq8hvYpN6dzfYd1B4jJ6n5p36NqG8ZlcyFTu
lhANlb09c4tKKDRuL7YSZyi3HywXVL3pAdlX1FN0KsJ91vcJBKe/oX6J6Jcy23Lh+eUOTSwxluDF
xG8zcSXxb7LSuutayoVZyTCr3xK+AMEDfeypBeJQAMK42xv/p95rWmXnQTMHnbzoG7X+87HOC45B
FmfBFwgabCbINVIE8B9aJEQpHMPO61TBtcGKqIDEr9j/uTVq+cqdsGprEdB0MtfGBIwjiD3nU4+w
4HeCBQAIRCz06jLAdHpkH7XKKnScZ+ZJ1kUbE31F3IpHlO4IYADoprJvlODUDHKl1aALOtYzBLFE
NXBfPKDtlTe1k58BLHviIge3OPSLr74Z9ewrhqDhH3Z9OT3o4odlj7AVwTBaM81mfQfn8QkSbHyQ
wj7eH9SPaRntaxAjYrlndqLCdIm136X+xunu+At7PmxvulFavxm1WP/+mpTSA6QR7CwYWF1Yv8CX
gdUTCh+T5WhclojO3L6yW8VjCdyO4DADEzvu8CUj0vUNeOME73s481R3NdBFH0/uxk14z0hITYOw
VSb/R4+4LAm36AnpCpX/cVRrk7PtjFk7uPFLTfHPifOu0loFjhr5Qsdty+0feRXyyfo0TQNKA7P2
i3a5d2KrkmmtKzrluGIP2CGqI0HCjzOipL7OZvzYElPPwc32/8g4YCNr7TFmx5/TfmJPnqUzoJxI
kB0wISYrxJFtfNDBEtUOa7T9pdWqDmfqWn2Uc/adntcp5HMPnp11Coh/TJyg7TsID6PZ3rWW5aoR
68roeAdov2+bdWgGIuy8keueqtQTRtzcYQk72o38QJEDsh+Gb2gumGzcyGvGOaFq/eBZj2S2hS4O
ts0meCNMeXZjs+vEPjaNjW4jIVN7o6GNaEEP5q8ZoQi3UJ4Hiq3ptuP1/oseIcoqTviQz+fCnvYn
dKzs0wTQ6YF5/H2h3hu5ew4ar5YNMzZWpaRUP1eD4MyGIHz0DEfDUPgCrGNx4epz/RT7t1AMoEtd
i/+5J/51MPn98UkFWHe2FlA/ZFYyJKN4uE4Q6sMRaE7Axi66Ma4oWVoasn+GwuyKRjO0Qa+htLwo
nsX3939PsyBI3nN7wsK2SsI7ckNZHukKF4AoPbmqOknsOqQAM7YGCAIjyWEftH/yZZaFEsDHXMfJ
PlS6viCzODx+ftWcTwwoOsOnyWN6RL2qpXmTCvY8qCjRHMhVuHKjs1+4v5orHEixY8zed/XTHJwk
XisgTLMMT0JG3hl47unXm3UMLtA7Mu570pv9stS/03zJYuV8yONa1elOwjjnCW8j/vu7nTmuaB7Y
m/06/bf6ryAZh25wlhoFCwlYSMne0UBdbhS1Ut/v9BHgYdeVEFojn1oN5VR6TjZ7lyVneMSlWAYl
n3P8kvpL/86coWGob4A8StYHGC9644UyAjqYXV13TZPdCS11JRHygiOTL+ABLM4pv3K/IrGhWc3h
gqALpIQ+4+vh4ZJA3KhBqVFs5ZwCtLvwAbuQhrsowASVyy4m6ztQA0+3hyXEL1IeaYFiCKiWmMBX
NFBg3gPFVFSMMy1BEl7xGERtaOAEmHyQ8FhKI5wx7Y20rnUvmE8v73RyCpMfOgmXrHgTIOfd5R/9
YW4OGbI1CeEpnvVTQ/0IZ3WS57U9UK7CeTez6kEaugK19380kARjjIl2tgkkZU0qCOPaZMv7NRoj
u7zuGHuA9WOQKSrGphKm1zwFeWBgVvdk8qvlCsKkyERsWcbpXott7x6NanLuo2Wa/YYoopbPhim9
MFTMrGQOvlYQ4s0qsLbaCfE8LN93FfrYyMoIf+AsNKjMsyM8jyLVCqsO9o1sKTQ61AP6hyXCQ7S5
BsUIMEadPyUN416gp3Cs2126BwQx239lnM43Am1MpAuionUbXvXofPb6RPRaTIbcvPDGhbRgFLHd
EsPXz0EU6ak240XVvezd5AOXmYDMLSNBzSBmEojL+dh8XRhx4b5byOjV2F+517vqjQ9o61mKxocJ
yHp4l6dV9WdoPZTakcMCiI8E8XqbhilJWfBsS9y09EOmh/3ItUzl96ktgO62c06+Bgp0mdppxPwm
Fh6XK5j1oaPWTB3+g3aF2tZOGA6KMT0sejWqqavMIBPd70LVIbspJSoSKyx5KpA+hmni8wvLz/3L
RjbutZhlwt6SNbVg0CMirO6iEP4G/lZIn5c38jD5rQ2YJhHg1Yo0yr4StfaryLyZ+JVyREDQgEHe
bhWdm41qT+V7PDsOCeSld09KOkgSePfUF0IohmJ/Wsw68VyQZcEwAJ2WK49RPC99z9p0bMNzdFVK
FAoiPnDyMpa1QxUYM9ypVit9z7Y6aZ0Tl0RCg+1losdtBG48V4Yo4VphxgIGrRCo3uQa5d8pIRIe
8oCSWLsmvo6BbTqWABkRpFCBl9I5zbYaNJyYLRpfS7xzAn8zgKjPAeitobhKbMoaUoe1lUfpireX
JKadc31FlHXWJCkazMu/TfNtOC0x3MSXqJ+/BAu+scwVHp2a9ofDQLlN3lecSD0wVtOLh3lvGWTk
N+7ad0CosukbTFzzMlw7nu+0x85cU76OlL4MJ/b3QvrrWsnuVTTQeKFd84ccuVT+tVW5Ra4SlfCn
ffEIKSCuzbOT/JR1Q3XSg/dE6LraRijRP1HcKhNvR5swBDeoQe9dHPq8onMrhFIwaozWhEQBonaW
vcVhpzabvjCSEX/JPthAEXdQhtPUG6D600A8N1Rm8D9JCBoiTdvOZbZrdAqi1STvTMbOGMDUzgCn
YaXnaD9gBcDe6/eJHqhnbyuIGw+5n3xCSRyrrvtf366KY6EaswbXkqGEXj5cc+FAVvRBGbGKcH+Z
HadX0GBvVmxQKN/pJvnEWCs7gnCOj6iCQVpJQhVZrxXu2UwYTxpEfWVRsP2jBW1G3Oh9EJb+5p4u
fA7kY8zweaNIN8n9Mzmd4BDjfEMEtUgef5197cF7FAUQ9ugI8Cl7FfSyTDiwuRDIJ+Td/YbdX1He
s+E23BUDh2swmETYeWxoglX1gKHOXmITk4JSnlwiKqGHOmc2+bo1lnpIkfWZgRG5wjUJuGbF3V6u
REa+T2PbUiLTk636T+b4wxhLV2vAbUxL2UVZxaXxfFwD+egvT4Akl17ACPMaQdAQyNfx5xFvq6+1
5hHZ7giM6qNVrBoc0dOLuqL0Zlod3lHpEgD+O3LzgrZCSI/5BzHcccN4TyBr4EhwdDOJfc4Zz9vo
CbDJq4aVzSuuvsYATzMtk0d6eNzQ/uQl8DAydcKGlHeT83VhJGmz7Yj3B7EmhoLzev3PxsD9Z8i0
YIpj7hVFrcaZgaA8Bx5f05AovtQZhzXwEq2qNmAlY4G8VrQiwm0avCa5BCvpEgBSlPr2k0L0nObY
20T1mDryz8v3ZzPEpbYQSjNvzCCJfUk0iTXd24YvZm0AEn/NkDfGzuLJVRDJwlGPgHTtlzmHn1aS
CHku8BcddE+cM7HiQCxHaloy3/mhOj1xHOyQ42OFrUKTI/FSzODr38zhYdVeEz40faLU5o5N7Cow
pCqyqKXu8m5IQf+0liPWSPnBYUoQ5Q2tVUVVgnVhQy/rW2Zj0YeIS3SXasKqOwPynLbhqEXIb7vt
q61wt6Cw0rNpDBmZTiGjwGNqBspvJ1MbP9Fa85chmLrPPv/WWLtz5Z7cYHYmY+YFKC6HhxFDj0Bd
kmqQb5cny1vszg6EsVLquOmHtE+I8Zg/HVdUB1c0X5wuyzkAaaDMsiMcIwye6dVE3/nNIc1m8VLI
dn4a8FPuNuzKXoOqwoVc78yC2gG0WnJvYdavzL49XWhXZziQPmfxjsxHB1KX8tb2tsh7vGv8UveD
+SFyjK/tW6qL0y/reWyTtOP0quSv9W0m2n7HR0NxfZUktgMOKM+mJQtVKf+R4TJHpqc7C568HBIA
MmugdWIfpQ7wrYWqsTwRlPfSjjnNM39u+k44Wqjcrpxh3BIUZCAyM6ItXM/htJd2rhJXJa+UaLjn
oEh6RogqhXbJ10QcGS543Ddp1saJNT63jj8U5nYJiI+JTu3O3JgMt2qQt+do+VN74PPkEUvQJZ/f
ii5UpGMEPbxV7AWGZgknytSeE/OG7XYOdaF0lHNOhK37FTGVDvFJ2/uyUcFOY71he5UaecW5tOm3
EUMoWCM+83yay6B/TNN2AESEZazHfd2zyXDWxr5sqgLFDXqzOA96TzMhiXvdmUse9kL9z3uWWCrv
CJQnheSjhL6j00SKlhHYlTfdncgTwjspWjFUGLjubWuiZd7JYwEiPw/Ji/vtsNyhl8uT1xXEaiCi
6LhzFIg415qMm6B4fM9gwsgyhqfw2QfXhJshN+MZBWoGMKuqNV8xJhpr2CKQRhe49rL8Eo3ztQxB
gMUZsPhle8pOd85S4f7lVa6ZslMHc+RoEPovIjBZTCOaH76Ysij7dR99FOEfM6GRKWyLg7EAmNiz
I4jWcxr7/fFoxNE4T4BggzXv7GIqqley8jDipsFg0zVhDraUOFfoZR+c86xFv2bynKjqLD7D/CcY
mbahYa6ZAiPPP1xGXdSlq0pR49s+VyujaEuu20N3W1gLUcPsRE82++Os6wc1mcinix2WnzF5D1P1
f7DUDayRAXEo3CYPfwIpHNkdPdxXKinH3FkoeOGAWpHGngIL8Ers5gfZY3NK+pINHv03Z7wctRL3
diY2P4rkhxqLPgvWaIm5XL6gUO+dNP/P1BbnLcbFvmvgck2gBym/oLpPQ/lmy/6RZHsZ4XtdpCuA
JgHp/7QXDAqunpERBHiEWJKFyfRI9zmmdbucGdWEmExEZLJiGnsqtY8CXJn+QWEgQqCKB8SR+B4Q
CdvdCNTd8KeDvsCpKqE2vLXCFyKuZrnP6OKlXaA4legH0VUutAsuOcn6JNJPD5TxZ9Fo61jhL0c5
4emXhR0Tl5MBsPr143oGeV4y7F8JeN94WTraBS710dMHuvHRrReJGk0sBYsDlBEHV6DGHbNNhTMd
iZaPezbiS/ll/4AqflQVC0uUwYEfgV/Rn52nhkoIpLBdWl5dqXfjg0FU5brewGqaMRooT7nXdb9C
HEyIngmXgovFzJYyUe7hejMaa/4lc0SE877uUm6FbpYlJbC8s0wGsgnLVv6ATFYCkhjQp43UOkMl
XKnINoTUlr6c0vB9at62IF5qULikdHacauz5VHpfblRDFwNA00VpxRwALDVytAwKjeKXjgaybB85
jAA23AQUSRUrAU5L9GfW0hMA/t6Ksnz5HIxDR0/oN+d7YqYu1CeT5gU2MU9Dd1eN8q5hrWBnRcch
cz+OZHr3Rjag00UTctG0LS0T1vNAwLCtnrjB4ICa824kJjyCFcwQTSS0o+XFdHg+Z6/9yWPOBkJb
e+cNdNxpggkJsX+6VkwcuxaplKW1wRYCoGhMe91NA5ShMdjvWwu2oRvx2NZgSIRuRW9Cb5tzyJ5e
S2xK9T7qq522DbRujE49gLw//SvOlcOILtfBAKoTkNchidUN2MSg55Q5Y/6csV5QwgXV9cuu+4Zl
Gq29TDxidfO/caEmtJ+ok20uRnjTe0hOpVbp7jH7YejUz14VlkG95tp+82NOwp6q46bJsYHf7f5u
FvaeRt8FM9SXxdiF+THwiaJARsL5Zru1FiTN8tMoRM2qGE8Lp46jXEwvX6TTRe5sSkzVJ6N/ecHQ
zHnHafP1hmXhEEe1tFBMyM3rSbY9CLhNh7keamzYn44TAPyrEZAkyOAa38tGfUCYtNu2sk1EzNRM
GDqNhwIClhKn9SbURGGbjHu59Unt3cHut1uq3qC69Mm+4Ia17LEZzkrU9M+Tj2L03wGz8JgwDRmX
neKb23nZvdXIQ2q5Gb5BTIvxZfaMYiXjRXK+WSea64ACOm2ezXVuLGMJZdeufwXbve59CUuzpt5U
KU/8zEgk9iogEHPaEd70/bm9HJh9DZ90Nos0U+YZS4GN6lvNN/3C+I6zK9z1O4VuAPcbZ+We2ZDr
SoGghC+X+tj7DDQ6Ga03ZVrQzvHRHqXxAQ+rb7mW7BYfFJ+FixkxkxZJhp8yNHOAC0TbL23q0WED
XfEdVvU1pAphS6V8/WJwh/K6ah5ldW7BFFkrRZ4+gh4RommKHc6LBpKL3S98kum+iAuNVM2cTl2J
iTQzHFCAuipU/5IgQ7CA9RFQmT4dfWTCzMfKlcZW3mcaEG4MHGMt3M8EHCAc9Q4rtmZFNLfxp+ZG
DCgZtEEOF9fhrvurcwWEEZ/9m5FHxvZLLRsu7bMaBqA7Z6ZLiMY2ZvelFdjS0dSH3sS5IYube+4F
kr6F+NxtOiaygI75DhGal3pw3tt4oVMzpkrK/eTOmlh6m7Ooe1aYbSJnQCuA/J8p6GHJe5fa8j6X
QicbA2OpnyI2uPirq963ovT9ESoeva59AunSg97R9171WhnTxf38tCEUu2BzZ6SvYd3tlSzWmxV8
xIqNUJNtR+2JvAcDfTocFy43RoIgxkBRBCILjQYDMxmPeq8w6pzSw19KP/CYpYOOFXm2/M1a3jqJ
S+Rzc6R/eCvIg2a1worQjso2CI3PQeIvdAzsI23JxlDz12GGHKV8OqdJBGXlB7SnyVy16SY4iIPW
wDLRSuXtj7Yk/1rqX/ZVL4z/A+RV3MY9E5Gy7jwhxN+JOxT9M8bRbxNhlK6Z9OWAfKkYi0ew2XPo
iMI9GAm+iMdP8ZpF+CoMYIl2YOS+OdIC1FwyGJ4h64BRf4bAwK+V2wqy8KB13kE2xdQGZLWor0DT
6QMoTAIQ+9E8vGmR9s/n8Z6E9gVSjVwmhoz8einMOYyL5uTX+5+eYAeJB6hydaVP+Lk/swj8aWco
z7UMS06C6ZKeUFcieGOWUCkSuiaK/Nzs23WrrsYxvA5IlI7EAkkSMKQhsL39GsynL981QE57XEQk
33jJVNaT7APGpW0850WSBls944VoJu7WQHrIQrWDtO1r1X8fMI+bbx/nMLvfgVTNwU+q/kV6ElWk
FIjf3uuwJG7T3ZGE9rkbLDK8yF06L9bpOS1ivbQqfRtlSc9XVDDoTBL5ijBOdc2SH2f64+ua/Y9S
8C0n8B7F2ToNHTFqArEmREFztlMq0udp0H6443URYd4kbtbB//Qfdfo5uym9T7skplRbHgbvXKct
H68qKvDTljQ4v5UVcDS1QHewuAVis6ZXTgUWLa2RKPzSe0StRfQ/zp8+e1Yrdu/xDiFn23vyE++O
ZrNLlDdYIQOuG3VAeUopOSOOInLKUKTqG4Ihj84wFBc6QeElFDF10VNTw0fvrh5Z8F/iiAq2onu5
/sZJhcC9H56o70D/T6CjgEUnXOdaiGKQUwg388cFp+VRSWEVHauDkQShyNl+x0DSwHqlCqbmpAJv
9yBj2Zoa+L9phWx1Bupv55ecyXCPRIYrcSoWUvjf6EfdIyQf3iTam4i75+/x+rIxKhb6a3P9PDfi
2lc6QnW6bC1RecFGMT8JAuLxK8C/4Fj/bRawQQ/CB3j66+RFjCY3QCEce9mUiCwjGsSILaXWRq/6
pfh3ftdc9Of28gczdTrIq9AJB7dbZpBJJAwuccvFtC7S48+FHOVEWvkymf4gBZEcpfaseTnonh1i
zBy1B2lK2j57MV+n9dSqEkUKV3kSgJOOfYIG2NnBS2lXVpa+2w5donA+uFLgayj+9EyHWLXc8GZa
DzzYRrteF2i/s5gnkb2qDKkoFzoCLBcJzw7ZBXJemmsT/wfDVLNxgW+3Y+poPiiwxhVEhFZeWzEr
whvhVCUdxASIRLUgobr4pBr7KJa+//k+DMnU7XYxtmOXMw1p9wpw2D9rvKYoEZXv6GrKwdUOcfJZ
c0KkBq38vIyA8v0S+ODDMbBlEHo7o8BHkoV7QVqI3hjRTzHDDv8qULuXMaThIAyfcZj0tEnIi7JY
FTUtFjqBVwLp0N0bY99Ay9e12UXyYLA4K7W5o4IC7YmF2yJgUGc3bOOPLtZdcAkhjTl3Wbx39twb
CRsV4BKDCTEDvy00cWuQibZHosJsS7ZW0C4xExsgLz8Ctowy1ojan4gIjx/PUfcf4IS2YMdTPUYy
PFlAq++CLaItgqGcmIUkmIepiqqUiWy8W2fvybBVI8B6St0MFM0DVq8RQeUfZMyaioasyCiH23db
KdRFGYFGoccDxoAPFWN44oYcAyylACoCO5epnqFLtc+VnVpPkShMemrFqbnrp1Z2DT+Y6zbsfmSq
Ne3+KyUZkaxe2GQDk8kUztKEK5PZ33xS0B+SpeTbAkoqJAgTmbj60JDT+5FGcQUdr3etpBHXJBpH
Y0yJWJh7Gybkv6BKDM2uVIpuMoAVmGS9x7cXYMfHOtoQdVGWwNTFo7H/Ec7aiQlNBPe3ZLu2JJUR
rhSpRs0jqvqmgde6WeLIwHVG8f7Z4sY22cvMsIxz3w9wL/pxusoCtERbssJuFnIr9BHej+kJljMq
mU1nwPMatHaQoOgEAuL9uzrWznxV+lCefqBdyOzg40uT7ng9lRcx3SKGc9eLHIGClvXe8/u4n5Ic
lgkM8VDKHGwmT0AaQ/yO1mwWDE+pNNRW+ZxJ5/kXks3mLx3yAQFpSAHjYYsuMW5nIVb5FlGcsTAH
teKKhO/f1D3WSHKZbAtiVQXGlHTVOiumnNYMNA+TCqQE32uKLzACJu7cHFG91mIGcmHVdRKCq+lA
NMN5jz19hkJY5cP4bcuVJVgXFmoyArJHKsgbrrRfr6vKtIvzWtJ7pZHZGuIg+H8aJgDpwWpbpGXN
+9OBHV/CVKzcLMQKZYv9NLJWKoJFjU2NHUbCBVVhlxm+9rMHalkygV0q8Fb7S2sm+ibsiajbSpIY
TgRIGwl2JDn7qZn/v1FkYqcFQsF4FRS2iM3ggdZJJlQV/16z2y+JdPSJq/Gr0h4e5P5sninO8Po9
bcY/mGGCSoU+Ep/V5pF5BzfLxH4CqcivkYTOgvtJZwGeQTCBlSk3eZtVkvkTuqz4w1DGAw6D3GN2
FZDo4exv/AkbXeP3vfK8mhF89a/HRDLDitAMkJGCw6nRMlF50Q+ItpIck5bRw8MDG17mTHjbpFGV
GT4fDn1uOwLLDJFZhS0x/Azj6OD6L4bqO8/fKy1jPB8KoyQdhfNj33h3J4ZX12w+JixLB+IY9qto
DK01azRGIxgjLHtsnRqckjJC14maLxZUScIVSd3dN+fN3BvhlDrkajRxTI27knQabhjhL7+r7eSI
TOGG1b0GPOLHKPTtwD+uvnRQEGz/Mu4NLE5Zdk4ZOoSZO4T6KbdBF0ukF9HbnyR4nICXSVwOYPsN
q8d0kfdD6eeamHb7A+9jRJPVvr1XG3rGC6WrqP5JARL4Sj9bkg7744M4afpIcqMvGcKqEtzTGv1X
UQOqSYj0CgBT3HCbqcW0w8T+vQmi0uO29xV2u0E1zjE3nzNbaxrVfinL9XgNYywcDf3jyd2I6AqQ
cVi39ZRKdNd6p0Y0dZPsW1kyGcMF41MDQhIABtwX/Er5M8nbK1K4ZWY9ur90C5ehA1tdQ82K3wIl
tyOIxx0GDThmb6e/AJaWnnjmLKk/ERL5WKPhmzxwtdk0md1Gk3DwZWekIPYhAVCoRu5zFnLhqNqb
xs5OStJf9NxzxXMPj7uosMSYCHi0COGjgcpA3lhQ+rgzXYb08HDUzVHkslk5/koLVY1rhiTAKLd8
O3iwC2nwIfdbTHDYnTxeR1PMqLrfQeimc8F0k/LW+aduDhWoX8/CjzC7NB3AoQmkcA6KZsZqnraJ
PvYBym7Y1CUFXYElKtfMFnBOivsE+hZPE5pmwgbaqFQ54XYQ+xmFkcbiMV8dlktmm5EsvFtdwt1W
ytHATSWBj1IP+FxjVLfBcl7xngrEU24ji4z2DIoEWu5k/GMJ8plGJ6uTPMcySx3axOl77G17f3kT
Qf95+6ZXwHb1AchJlOphSAhqkOTuQW9Tp3AbEuJ+61qldw3FTaJ1woudwNcn2X31dBLOnIpEZRFl
O0ZBE8cysuXaKpUIwB7bWeR33gI2ac31ZdBGuyPZbFJ3ElRgusS128b2dYaCJHQZIxKqYkOAFovW
LpuLhgiFkz5TLDnpc8Bl/xP11sQNQP3nvqvA3HQtwJOn4cxWT4tNgKZdiZ94UTE9NitxtqyGGAVU
VTP4aBXyNrorrthasxeMKkQ8VT2SoVGuc2J1iYrLlpyL1pKnofq8Xsl/K8cdxH/Ij6KIUc0hMpyp
DxviqWmqT567fPXxIJmSSSEyAv1ydxc2mSZx5pbZuautubtxXsPwikeiSiDY/dJnEAmR1PF8pSnE
05re0X9dCklxc5JujIxWI//mv5CXSLYTIM0+z7OVliS7xY/XHhjTY05DDogvXwycM0lWIRQETRNm
XBB/l9AcClJfosvxdYzLZmO0GMAbHoz4IOIUiHvxSu1vXetOGmiYFSEl1+fE9SqotL8hfX1Am8Io
zNikBVHNnRzsOv0Gg0wSRRJXbSKdIsRu6LSB4+moofBy/QF3rHOcchRSU/mk6DXt3IfVh1tJGU56
mHWB/ItQ+4mKmgOM2WLzqeYX3lfSNsLhLZmc8tqOrN9/OZv/QOG6QjCqTE1yYdvAPz5sKYolZ+bS
w+aMzoDg5VD+MvnTxUFOY86hYVDKForob11HBx8iWgQZ1t8RRVAMUwGCyL+Er5JjmtxbuyyT3H4I
nqGLzZXyqZ4TQRgk/JXJQ0O9acdarqXca77j2wtJlta3y1Dv4BHcp/3h2MYrItLSzvkg2jdL/ZwL
228LsbpKiLHCws+pQfG6tKa0OqDqFl+HQXrwCL7YUzOA1aqA/SYA54wG1CPgQ0lT/M1MpL60emkI
ysXMpWPHCHFUjpS0INm+FCJhl84nkSgFESzDI5ZKJeVzkacpk8zJxFzyKWkqYZl50b/xoeOQZg31
5K8vd9W/b/RMYLjJCzc1eFY6UQ9oe8hMm0rvUIOtsWd1dtxPAlMFEfpuul8ZkMCLDas14iDGZlHe
jo55ySrTczuERwYR5Bb/028XLsFbzYXCsalE3xHLC7ArRR7AbYfZdKlzoBLVP/r5Ckb+kOPw34ZU
v6LNuVDg4ESdREs5OkXBueNv8TmoTtDh/wys2gYbilFOSJjHam2bKWANFVpCpTmA8+mWsJq39akb
L5CSW1KGLGzF8rI+UPyjH4+g6clcVw30chsV2KRkiiBVn5H5kwI9+hpUteuUV1X3u3YS7CWahC6t
/P5h3Pi4v+F0fB7Qj9abL9gAbWrqS38Rd9JdzCODEgyJIiwXmlKAe5M/1MRm2aIijQ0mVk3FOsP/
Ur93vTmUtvX0XUdPn7Wh39DvgZKMEtSw/UkhBaa56w7d4ug9LraYTmAszb58CUD7k4hdwTt6VbiF
bloRtbHvHkKQuo70I+q4OD2YYyFrfP9FUv7z7CJmLw4+WltASF7+abK3ARTlCGoeamGo2We+Q9Bh
+ByyMo0iSeqpeKAMdZ61kNZl/Ah/pGUI2iXfLHJDeEqPz/CcI+9Otf/9gUHbbcyfJQDkYHnFNah4
SoiF2wToJWDA0MtAg+bl5Kr0m41cgM97eo42QLSU359hy6lnlGBA7WeEli1x6AEO0bHZiqsCkICX
o/gtqKq179iD5ADM+u442UnLQFDYVuUuu8Cuced3FMShZxYh6Moel++1Ld7K7E0Jx3mfb9nTN2BM
mPgSDLLEpSWht0xrnppuJ4IAqVdjMtzm7mgbtQ9PiN/GnYXjJGzhBH6LTVsJw1D6W3U+F8vjRiZx
pJK3cfebUK5giFKstBPSdjrWeRAqoTG0e5g6jq4fvrfRk4r7nLJRcR7nBH4rHfMecBBzODY/n4AO
gjLgX/blheL7AAcvIzDr8//HRFSX+kiGi9PccLO8J6QUbnUXu9jeZ7l02Tkcxc6mc65eaA4GFdt5
mRTsHL/3XWmqzbedaApODgTOtGwsEQHUefcPdDPWe2OVQYnnE8WrrqjVMz+2h4rNnH/NZ0G9QKsH
b6HGYf2kRMLYXNbC5L8H1QHIlqqskEjP/i5rP4czZYrWTlgUjP2DQTOV1Vw0KoHSHuzv6fZfbEum
+Wz9j8GTBgiC6MiaWwS5QQwcu2KHYlG1uj/ihpZitssDP1vlCM+lMxpyqeMTG/HD4ulaQAQVGqxS
ZSJs9TKjiAQFUzVvrziJ4y2NUMLy1uA0UuCIq49hnTy4mpRk5WOeOWJXlm+jkNjQZiKoLWWEllEB
Mn3baMq5AY56D55oMgyPfYHpS09IWPdBHwS8zDfY08/AOyvzz2vHh5sTxh/l7V45GbqeZN0slwby
MkMsoPMINX2V8ndLxdKInYIv+e1gJsdyByu2pghdxndnGt/AcZGa9ZV2HVbhCbyUKnyFyNY/tn4a
hV0eEpY7stZ5GVYqHUUaM8qqUhLwQp8M34ULTNJYomFIOufrGIg91LInbnNRY3tlsFGX3dPYN7el
vqFWOpXqKK37Zy5swY55yTqKSdGyVF8etOjZE5cXo9HR2FzkVogMKuc3Gl48cFj2vK/WJtm/6mLj
LViyQ8MtocldUjZedw9J/QFxAFhoI/bMwHsK9GmfU/GRZKrlK6hMmQwbIzNk0j75uToQflQSSulW
3qQSvuXRTn3wSikz0SkUWzp/fnR80Nostsv5LQVBgiEE3Zx1Xs64KCvPKfJxVAurpptPh8zrfTOX
Rqf1U2/oanYFnIp3FbWbeqyk1YS8jeSTTYN6kIj3X075ZaGV/2+rCWQsfFR7u3Q9I6gunwzQfn2b
qQPxt/Zl48c7v7w3nkYg1YfMslCPQ1YeZsqVLo8yWzsNV4WanWqytFvR+uLoHa+gike0YVCmXG4a
J29wkAf+HpX2RiOS/LMHUz8El4ylI6bzi+9HzkiLlyquMZVTOUCF5mNJqdN/AgHJgGvqrxFbK5YO
HKLg6lBrVy8MV9ueWn45AHG1RbI/Dp5FS+sSbPiJW/hqiL7e/wMYF4UvWVfaOBbOcPlK/spsc9sq
p+wJ9/MwxTKdYXrpR4bEOsWsu4LA7246vUk6Qf1AV0Camoey0oeTjWggE45JUNnpt8NkFE0yjZjq
g9/+xlakNFs6v7jBdGl7vk3o1ybgdGpmpPJpJ5hFaapgtLO2ct2cJKs9h28PAWovJl9kX11qmtDA
8g06U0E3fLJNSOdLuN+7UGGQkwIbR6hQZO27oAI4YIOkei0jzA2h8oSfOImr137quwtG1k/Q8+T2
eaqfl6JJvPtIfO8M4O01zdNfjTtdeGDWCyQpHXy+kjnSrFLVf1W3YQsOph+e2xbH0LuzlfaLgELj
U3g6m6Pgd+9gcT8FFFEfL8NYmt0TmqZjHROgocywvjE2agOKh37+PHdNhzRH26ZUmS66iYVU35+V
yfaoe9LtXz0n+FjepWhN0SksQRVJCR/CXEktaj1sePoJYB5ppttcZ1VUbvFbjDhrfbWvqpW76Puw
/kmRWGQl0OFAGUh+omQ9iLpMFyKRwYuStPIgUIRSeVbhKEFEUIaMSQrHFSLCIML0cKOW+FwSYEzz
mLzvpzZE3eZcnvk6HuyW2NMZGUYpHpMCI3FhbwG9U7/hOWucEj6kMrzU9wnNsD7VV1L2TfU6TG9J
SHH6LGyijfAW0XonDNqwq6I/8xk5q/R3AgRTmyzfyyfix092b9NutJy+4MkUfZZtw8RUQOikZjVZ
9oZ41hBnmgrfGjfoQ4rJ1g9yMbS37WaKRy5X0cNFL1yLvmVhejN0AGY5GIjT2RTo4UAwBqQuXcQt
UAS+O9X2fAdYtrc7b8v0rwqyDQOFi95M7kHMvbFgTcUJgUbvM9TnA4sF4VGgtpSNqL+VYovD7JSp
xGYF4OMgE0ukvL3E17/nQZfijfvXwlutfRlCh7I57nTq9M4XMry3H9O05WMIucRpGWo15IDNYOn0
3FJ/Kq5YfaLWAYDKpxQhuV0+nr0uH5QzM9Oeo4Wvr6AhvWw1SvTcA9QA6f2hHccK3EHC6leCj2Ij
H98W4FXmV8PXQMM3qnj1y3tR4qiAVDIDtJZPboemzacgwUy0RhaZcjcNV5kbGOgJNFwJdlZBQM28
OPuennizJ6O/lzcXqqiTvzca+E9bYNc1FsHwB4dBmvvj7VKVLxBn6OnaXWJr+ZeEATu5w2To/qWB
tl7cef2Eq6o9Y323z31ur+UTEG5Hnm2xKn+N1CEFCLeyy98M+d/enG7HszGPSQB/eC8lcsWZ30V6
0LfDBGz22Z8PkueSZzt+zWC66qnycuCyZPIVDJZyK2ulpqiSuyCamKlB5704OwM0T4AZ0GWtc0l4
y7QABAzr0oVlz4u6h8JRBA60vXO1VEpFH3obQNtcrilgftGnByTqkAmYuW6TmUhHqh9geXNIE25o
NEEtZBGgeNQC5HR/gM0pfy+gfBoh7hFaJQFDMhyAcqeKaXomT/HimWEGGLtVJDihcaDCbEuSlQos
YtaCDPqgZ3Vf17JxhcMuE/fFotnDNUTNkAJBQlNdzOt+Ia45aQxJ0E5EJPRAFQoog8YU/+qMCP93
D3m1HZfiixXFQ2WiGVfne9Fy6E120kVE/Gx3gEVWAqFt60GIVc9jFARLOWKZnYKt9128QmZERHQm
a1t6mO3l0MyktEeB9iUccX3jBMxTRrbbNN+IA7E6SwXyjjloRfp/hoAhIJdmTooHt0WWDEgAe/ve
jUl019vMr0JQmoFES/q02yGrYmUkfhw6Ls1EmdI4V/epEXgDPrS7SpUGypMy36JGZQs+KGFVpKeC
8qx6x2hjsa+sz77KrgphnKRgnGxNqtFaNqsbHffkWS4Sl+hxy7BxGmQQ2TETLXhEeF1KNHHjqlUX
l2tRMmo++YGueG7lum1BImYI+LEdrdIlVMOtq0UsW3aAynmTCCSdtRUS/UK36HCc4A3DcgoLB62t
lClMDd9zQkobXeDBwgANl3XA7bseuU3iyMXSN7dPdNTIgk0p4fbSUoyz7y+DbewlNFwftHi6Cc/Q
KATxSsCoxk3zBf+7obQaD+cXFHXRJwADiOvilv0k9i/6aOadva/+0JTOecNQbenjJiAXLl3Vl5Ov
2wbWfYi7w8ysIHzTphMYWzWB3PGcVVszR+1zYfK1UazkrJcdTCEFz4tjehooyHXC8EaM00M6HVhj
+89yPV24sMekDU9Zw1aN3YGDp9PB+8mgg7bzFazvknfuNpTs4qI6f2Eukour/yV9wG/7hMzhBayQ
aEUuEkAkHswpRNVp31C+uyzwRuoGUodPGUXY6kGU+W/RV9vp4j/gz1TZSz3gqdFDbE/gqc5kS26O
4Np6zbGkMYJ4WjsE1J4JtOElHja6DuxbMvBmkOjWhs9eGfwcvgugJx6J45Wu8RlAT8qVDcGVtgBy
f8SfKbPw22yGBtEGGBajS8mCGzC1sRhbDn4RKOKBb8FiBiDZrLoFh5vOJVieIHG6lGhz//pTqvHS
DzXUreOKeRaiX6aAJanj00E9/NLIosZbuJobEGqBG5L0wO1uYxNm0IR1lnmhU71bg2Mbs2SWVwR6
RMlYGCxPslGc3mRhuo4WUovOFtjRzomncftYA4IwTgMsonnVm+P/S1FyIFGQuIuOJ0RYcqWLnaxp
oh+yNIgRJykSwQHbp2T/IfrNJZo8Sl0FYCG5UIFEnpHCH2NOpO+04uN4u/ASkqqh8WONSEwpll0i
uUcX6AvnjEEGnl82ll2py5qT+2F1F+TSLuS2GTgBmlxUXVK+lFFbajYkXXNQWckN0DN9c6/mPgZz
0+nZSKcCqlbdeGc7AlwiPapo/2UkQbwI1hUk6jBJoh2gseqYQMtKeOrey7FouduAYG7BtqTNIvbg
rx21m342PQA7kGJy0nybEzTX6o+W/+UaZXPQdcSs4xp+i0H5c6F4CBPy06YTjHT5V+O7Vq0XQRk7
ekbpfH3rQFABd5j0hA4N+LFwDbR8tUgbo+QUNw/gNCVx/8KwAaDQF/ydNk1C8Qezs2iWV+cOvcTc
E9UhI1vbhfPGTeZIrk4ayfTQh2Ktk28LazdcD3u1l+l7cIeKtjEkq6+N+z3/Em41QXUvDp77jGK3
WxC9RAyjFn9i8fmfy7zcCve+2ZkI77JST6o8Z4Q//4NKQ1mpTivvDcFDFlpnn+x4VTilGu3HrHrx
izgVJPZVJPkGPidXsIUZkS291dhf6V9sYhvYvSuC9MxbP1Sh8lyqvrmcbBLEOyw3EuiFK1X6y0VA
DHJOAyXYQLa+xwH7WnoOBakCsLo9oT3z6i5iSHfinQdgtHFk08qSG5dJz2jAppByQts8llSKhSOl
TheG2DEIwGMeia6PHZRr20POknFTmPItTPx7FB775L1Nc/AUFqRDqhhwNtSj3+ODFt/fvTmswPIg
u0w2+VTKU8cMSnSU0qLsisR4nLPkOdpjzZFa9PRnSMrBQHD1jzlYQFT+Qj50PyIjQbqesxyphTwR
tmUXwI97xkU7I7rXLt65dtDSxnqLVymMBKH0FkFLwPu7Ecc+p8X8vOKx99e4+A8x+3ZNqDBMRi/h
JWTky9f8pwdvOZZEufw6y4zJSdZjNixECG/53Acv6kEsAmrXj8uwi7smdeIb+90WZQse1FUTh2de
w8Um6l9Af4Y9l7+lDOJeiKTqHubeam9IXsnKUjPU0Qo2cgRxPWvmSCm4tCjeMTcCWYE3bi302ziI
xrsgV5RoQ/rDg0XkraGMOWhsBawvM0ayudpZg4NU2IpvcH7wMbDollm1f8AGxRY9gOHvNWoyt6jK
ymTMtTV2p6UurbXUgC9re+iAbT4RQ1n2VNKHjLmFNXL3PvSt6+iEsxZXhx397+ixVvP+3E3qsSqE
JpLukGmdOojoLp460zf9bWUsHjXPCvdKedkc79+EnfqLzMbyEQZG05O4SNsQEQYNYyRNhlIL3aCK
JFGmWIzlj7n+xhIot2pDbCt+76HvlYJIfhksFpJxjC26dGGmYd6u5g7VeL7CWhE7RYPwZU/YC4ov
LTVunMNU7xEOONh3lUYlgp2pr1t7ISzr6lq8U/X6MCVcIryTaDz0cdGCNbXKyuYd1qjtY5kJcIBn
/Pf7Hf2I09trxEdPFWiJwR6byIFRQON/1ZnmfoxF4naD54e+emywkq7tX2AtAFAYKDXMR1Q4XaI7
vRC8tI65AVSbEvolx9qBysmTnU5JE72bZglVb3gCuBgbbCQkb77cFdLHTwBw5DTVTTUdttrZtPp3
gwAx+5xyT1BiD9Qe74zgvUZ4Fss+m0QbuPIUPXeDfXo1EnRDg2nlx2xOBqlU1QwOqw4aBgdXFcIp
PBTLvwlHRYxWPBDxc+bM7J5xqVfQBCp2OBlFUkuCuhuR1zwKRFVMgJSRd2TW/Wg41cndZnPmsC4L
oNJBKKtQFJXpeVVpoPbdagXAqIb3LNBJvzBhIADlu4ZTwGMZLfUuPXBbL93502dEML8gyJ/zxu+7
5jRVWkRohy6Jxyjnml2Gb4UNlPXVjJn0BzKwmisBmRc8QKzGMyTsyyCAu/Bxa1B/2lAMnK0FmKS8
RQTfmLmXrwvWQ1ENTrfQFqy3MvM/tJsL/C6begDyG1g433XM3pe1pYqQG6pXeI8yBTZmZkI7qq5B
weKbUqAKq7P6ujz/tTd1sRIt4QOdkUZ9FB+z6+rfzef3e8zs73s8XjVpr1SrwORBb1szrE1VVuyl
s8pLJ8gxXy9EOsKb8n9O0RYqxg0Ws+X9jWdqmgijIvKiWSKzB6jLPwtMvkGlqptiJD8LZ6ZAAlZM
PUgdjzuIiGAMoA4jhEpGcvMiN4LHEYHvSeWSJ+EQR0V84ovxyfW3Ot1ea9j3PfygX3Hzx6dCRpR3
o4g6AV9XMNsXbTuYZ2TqJsH5fPt8qm91tG+tdefc5uBP9Y3UEyoLPqQuy+gLbChU87/31gUy/6U/
yVS0mdkl/RYzdSW3j8DDhtZThvQCQx+S7HBK0KzfBMGsUsPvLgOUYIZ2tc5ZVXcctgCWJJE3whqG
cKkvE6tiBKhH5J244r8XxC0LQcOg4vs/h3Z9NkOhdvM8rvNrxEFJAuU1N0ymfUjiVmEvRgA20wWd
QTF0B8bSb7Kv23IyXTrDSjjDgHCw/9Hna9mjcLHezqLSSUyYSHaIhjnr5zwOopmcI7cV6Z+uJvqy
8205Dz21VoYNaNQtjbNWlznFWoATYWMiB3XIP7zGOTqzrqTy5rvsviPhawuVB3mVl2f8yYTcaWWO
ft3jddeu6XGX8B2N0T5xhl/catzxLrSubwIG44N3hEh+PjpqrZIOo/Nq0jqf5pc0UMY4rNPIlVny
/iLVc1Qf7dTO0pQ16IIwsZDi2sqOggOjcNKBR2wOIESD/W2WqKCzMDrCzk6Wb0zVVMG419OrpXwQ
5ryHNTFmSvlCVsENURxeraxDe/Fv5b4/L/dNpaOdco+helCZjdRfAMPbjU7KK+QNrzgLDse2qA0M
LRqXkk/4Kx2oRDmTDuQPMj/LN8HmhHzLjJuUErR7KckAFGGt6Oku4tVSlstdPHB9bjER/F4TozHp
D1I66SQhcxmj52737Rev0PTKyEKfr/Zp1nFOVJDspaPeOjbMGXtNzyd9PEf9oEbec9hqMJedux/g
Z22QZa+ufUYzv0w2Ng519rJiHmy9l3mhcPAbxCWEA/iAxrlMuW76NN50T72ZKntyP1dIJfnxtvZp
/ukxrZmkmeoQXeFVupuiYKxQqVAAqUhEAWudbGe0mmEUd3oHsy6cP4rOG3nGNyJrbA7Tb9mU30at
AAFFSBZWePU0430x2A5egh3nGvSojNUH6+h4E5Wd3Bao/ywZ+ytOyIEEzZr5qfsh1vvJ7LSaydau
IabhsBeKs+OVKr7AommaLU9JwKWTkeyhqHFAX2mgTLBjR8cZeAR1WbU/vXDIvzCQM+kMg/gNPBOq
DkhUi062ShuOJlRlK8Wf6UN0+1F6j3+sQZgMzxsQE6U8ZzvqIOmE0MmaiIUhlPvmUKGmcj6rS6SV
Eo8Roc2STzMZSvNyi3LoFN0faKbkky4C3J43RxAhpNATGtlU91bx4ZcnjLQEj/R4Ri04YC+Pv1JX
KsyzyoRTIkI1dkDxwV98VbGR4vMTrMXQvY2Si9I17bksAP4/FBf0+Gkx3zd9nd7YI8rCLaBSMTX5
NSc9ZHbhCGznszzOSU/vQyxvUyf1k1P7a/oJuCw+SiLCg3sEIHlh3kwuPw8YkvTZD6PI9OmRbT9q
w9R/AiN/cH2WfXQCA4iK9ZIqS2hJvVBoxhfqZOxqUarqVlZiwxEFa5Bmx/sIzVrE1R2tQnYhm1g6
9IV8yWTBOgmXW0g01A97TmufbN3d090Ju9E2gwO4X/NFRqXXQnvGbMXN0OcwjWwUT3V2vLM0tF3t
Dodhzrv6swyHNqlXXyWBbJTzYC4V92MhyhiGVVthI5g6IYDJKOi1Nm+hUR8Ni2swTHU+u4IGji3H
vE1c68n9CDLG0W5ksBCr6DIeFgav6bFeEGxU/9WLSKgWyZbXWBxsq4IuHEK74oKdbQ0fFMOeOtW7
/kPZBZuYNKEk36QE+Fw+0fb8FFYuft+yA2Q1wYTX832WNcZZmSE7VOyvEMFShawi4agMPflgmaAX
5zsaggFTew06pze3Hobpb1Lr874ZhK0y+sSGAs42YwBmtlkX7wccZmOW7Ti8cNMquraFnLaNMSxL
FY4FxGTcdVpMLHmCvZHIh6b3/J+qGN7TLXIgWcip1cY9Wn4BpFW3OKKyh9t2Ui7dlWsPoc3WeSXJ
zPGFC+2goclfmQq0SybxiyMMpH6SIBJkMbSvuUWq3I+Ckf7KD9q4NwZRrBgkbXkcEmRzCpLXo45q
fyqt0W5MxTofCZxwESBGdLCFgTKzX4vrgVSdbaflAesga9WxJDw7v5TEM9FkbaWIIM0I4O5xDfYX
fdDS7jA8JquHXaPtk5L3WO0MxDnYXcBd8Ld6TgC+1AqhQ0xi2se6W7y/I8Ca4q+dZWYqOAmBuVko
XHE4R4Xb1dfVhJkv9BkcFjheRBTIwx+ZsYAl5I8NUPcfoVaURSzXtRwp4JK4sfHO/1x0yhBHtWuL
roMH4rMwcLzayKmG2JMipT5qqSfz4K5MxeoQCyZ7/YD1x9INgz91kZQvml13F7Zbndbdd5VAdlZg
tSwKq6fnZ9rMnbEF3FNhJuzvop4yALuWVJtpbzH8Bf6Wv0mjxxWdACfSeJNWOulFLm4SP3vKLuLk
FaHxu6WulVm0HOYpe7jP815IOJIRDzEIQFVtIwDC9cv6DX08fNKGbe/PeYhQndP+AnEChg9WXMWh
RJUDdRRIsUTXBKiwZbrhljGio8b6fdIvQoVd9L0Ljmw6Baq1rDTlWHCiywHynkEBYiaJx9MRUg6a
vT3bC7rIY/j9J6YbRDNN2U8PNG/b7QhdaNY9qm/urdzG1nJTauE2qY4AA5jJnF6xIbNrI4HtThHk
J4bWEZLoaKhmYO4ZqDXotLE233VUkxGLFIAoT1SL5DNru2IuMsK3sIYgPU8hSbjfnmbVl6IuEiL6
459SShRyaMeycph1lzu9++AJn42sePNRRFmDGYt+D8QbJTGORoZyRtDy5c/3vwKJd8v4zeFMrJhD
SkQ6KLb3z9PBLGlEym0ymZk56dukPTMHAGQT9vfPRLblv5bmjiSuBS/8hpsWGKhPxGO4sKjUl0l8
2axslrPTgGhUqnfMbMy+E81mTyHLiUGXh6PG+CmGnjrA+mRx1k6mL+rCR5SsY8wqFLrM+lhscoVr
UbyOlZuGw1TCP3KiQHBn1FyBWfrFD4c+0KXC8ut8O3W6Mv7FuzncYubMV1xfRnFQ13jwIIpDBq6X
exJMXrP9lehlBB39LV7mDjh99s0eBwXBCnjhrPQth5uAi7qmZq8V68xNFoKoXAp7SY3vPriADGZE
nrpvZnrSvNUesShNTxoWdQYxGeD34LD19Ww0fdevx+szz4fCNpa8WRkKUb2vfxwB4IKI4yzweVu5
/qySNWLDk3kPq2T6V7CihwDONd9guU6qx1faTgpjA1rkAbtk7roU9qatbKKfngRL1MjUZA3By0A3
Fgze0v7x4H07y/kL8PLFWTrCP27k+pwvhi1uQjza2r2k72CZvYcCFqQZ/VqgKrmKSWwMRxcUTqwR
WlKRfaUrhZhqcc+ON5reF2LP7tJXEsi7Q/TKrUnZLlk87GwpFWEjVcnTJTQ0KOb0aYSNPjZdwPCo
wVAITwj3axTa0i+mdEhTMGhYzN9Ka3Y5iSRCK+wBcT05UWxUqEJTHMly/2sQI9Fqpud0lCoW5zRS
ViYd1joOowRlhFQINe8rJBc7ZfV9U9zUD4I9qp+XydSx7x4/yOekSl9Zj949pDLdeFHjmNV6BHnx
qCDtiPXKQkE9Qyr2Zt4yAKdeKT/8YaWjGEobwl2e9diRztMb/5WZmDtU19Jb9YsiGkyJeaWLXR6O
266x+VvPOcoArrpAUp/y2qUEEhL2yrCAqn4Ct7gPPqefyf1rmOT67H5DKOdbxVeGVE5NMIcyfDJg
a/oV4HZn80ixLG/xL4WSe1AHBoliy+0ttA/oPYrbIyanwRv0ufYUxotfz7Sj4A254AGYf1bEc6Ku
OCC7RtrQJI/xDb5jIswTjtRmJrejw25O1ciu+9UbQKmNrBnMfEzZ4V0KLqd3R88i7VeQK/pVjj5J
Au/D/YpsXT5QaoAE+e/yt83FKn+7B1zzLz9pBFhBfCKf/F+fXSOY+ZbpwiPkPNQZjE0Ql3ioRn2J
bkX73v4wSnHs+h2rdtGx2Hj/XRDTtGXLiK3NrWUZxw1ycelU1JMOF1I2qdbVCK7H0G1pRl+hO5C3
p+je946s+ZEuH5Ap0BynHlbr3fjaEWzjqbPKI0ELvk3cxcjJWrtz7v+uSjFpE0ItJC0Qkt2bh/M7
DTt7GMsdmLyB6HsiGKYkyLchQ4neHGai2PbQjNxeXeICpWMZ5prmIwlpnj93CawEIE6UYBmW2Pcn
bEW1K775GpAb+o1H43+KTz/eJqGuzMF1ssdBW/A8yM2wr3xi7NeXnCZC76eZYfDdluLFhvZLupWz
TU6+MR/bcTHAiJtdGlY3zzSzRnw3ckPPrhvc/XJxj00frkHGqhN22YRtCS3yOZPmTahwHZTBFzsE
SPz7P6b9HvrzAlHGF89nCjCcT0OThgKgUZe5MCuafA6ExlFYzzd0ksG4J0MXiSsp29cUcJLg1TdA
lR3yLvlOFwLgwwzzlXVv/dDwQE/JxfLq9GEwbH6ihquf8yDKYYtMF2JZFmAMIzLLtuNhizanQ+w9
rBOuGvIr9wpIomfRLyOv/crVJRxvG01kGl8EwgNw8eCqj0LR9/g84+45TFPYKS2gQn6uGmdwRkog
hkkd7Cv7qriq5/hCGb93RBSAb4xKbAM+5gxphpHM5cvUMSfIUs2xyVHI00y8UkvWB8BVy44Qvr37
vEpsYt8hpq4oJm8julh0DLj6NHnemEUiwUXaxh21hGx+cGlumuM1cHMf9SG7SqdkoBg6hDwT6DyJ
El0zILWZPa3BM8pm8pmjnNg+1+/8z8Z37k8ezHInls3/Ow2iI7Rz7TdAEst1IOs7wOuIqaBU5Ahi
nfTF8dkzYlladxTfXNZes8q33mLQy25Rq65qJEeVKbtzPuBOPvqMnN6bqoaUY+ZBT0EWr8TQWTqY
FJctXg+gKuxp89J5nB9Wa0aZLqq9I9tUF9YE2h4/yI3MPkT/ZqkUa4gC7fzZfAXgn6YUwtaO6mS3
A/nN6obxfCU4GQdOE6/i/Nf8JgaFtzhM2yyLkvceJDvjGgABk/EEsj3rVf2Bk5KMSPWQzT+4LvZB
8zAd4NBg4wYjLBf2LYPWiZvtiIM4WaO9CMFSRXG1db03Uf/G/RWC1tSfizcU48r+wFqSydkCEXum
/9ROMrzraYqfP1BCptYdhdFYYrRVR6qucjdPIlj+CwatglOAdI6CpaeuX+CUNeUDlLpNTI54lHxi
nQJ09DXdGI5lOGwEX7YZa9r3i/bB7YmURf9jTGdK5xHnNwAVRAfnlZBGgE4JrTJOLn5k/cpnDVR/
5VHBw9qApWbO/lagkH6BXgPvu0sgDl5vhk9VDcwoAP2+1r4JAvCLVkGXt4SVitBBLnS69O+7zxWL
dTbOXgDAODTpTJYqFa4cCvrTX/b303kIFQZxtN+s8WTK1LVIQtD4P0/qa7LN/G63lTo6AOoCStfz
pI7j19k/c8pDRHV1mk+ZcubzFmez5XtmDwJ+gNZlwLF5V3jWsHo6KhaMEhfT6dQVKKeucQbv9342
u0grxh0p/jWIXj414/bsEB9tyx3EktViHTJf4gqiQU1GOyNiDyuqFzM1v8aVeR5AxTG9AaglsYs+
/iraa8F7At7Cxh5X2iHE6FG6On+VexsfMXlmYgUEH6r2FKD/JOgiMY1uytUYku50xSvPt+a4915v
4pygrOtY2BG7GPRDT5iFaU5+jxxrZeab7pEILNAYerZPdYih6J3+9O6qDCCgbX0mrx6FksfUU+kq
2yXb1iaCkV1fpkVL1zglob4g2bby+mk0mcU7rWyyhOSFTW9GuTHSBGuq8YlTUloY+64JVhN7dzek
l19RBDhY1KROR9EEb9Xz6YgUYpVkwELUYgjeqrHCtC//E/Ssewj56ec06jFZXY9lBaBDRsHNIrav
iDzGGofusbyTXiLAMaEKcOw37Vi1cc61xtL/aITsnTgwyn69SRJEvf2aJZN5JvDeUTbW5QjeEJ+W
tixr+3AWmRVtRAY/+PNkMywxkqbhFUryWAin3saBEJ+TzgaraiYSsNrM3f1xpjrRLbY2TuPIWC2l
cIU8HLWgqE/dB1myj1Ghj8IIyiIYG8NauCdkBEhhj2u4r4ah/NR20sLocLYYIFBloSlqNgqcjnZl
PGCtRtkv2N5YscpeDly1lTiblAaXX51Y31+4o8Fos2iqARfmUC7HD6j4Pjm1A1sd0kIl8GKgxpGR
lGCrgeV+jTbDdlooVhSseLxtB7THF5FXYL29cHa7JCisCItkNbI2iNlP8RwPD7sj/G28kxSWusjd
1a1Tp2jO/hNXOofr3hCCwgI4Us+DVvDGYnkNDrDJzHML7Hjhc5+VOK4eRsAHMiwAYOI4t7Z+bM1v
iDzhYufe2GndK3soP803r1FxCZ1/PXg85qweWkpXMBqb30gJoz9ii07uWkn0qzY76Bffu3wx69AS
srgX/Up7sxgYX5ZsZjARE+XJL2BlSPyvCK5GcK+Hl5xvhG72BaB8ghNw3BN43VM56bKkCfGR1keK
cyPJ9uFlAnQpbZyBOeXmyg/TnxL1FQnoZsUOYNk1HI+Q6u7nzIbbFkmzaBteES63OXMg1Yd2+p9a
CsBDpkMSKA0ITVX8vqCG/psYqdxjq3PU4oF53L+1N6XYkok6tpe8SHQFw1a6mj9Bp+vy6fmMFNBw
MqrG8bxtPK8zMW/0uXC7AID+er5Aw37D7tpjzj0KwTa8X4zrcfzGlNe6V0KJkYMSnfyGmSkjoqpi
mJEgVzMlp+IBSK7eNj9a5CSxrA8Vd5A/0gbQAyjwRXmqvsxGOEcpcs+OBuVAfTVihzrRcUixXXyQ
pl0vlN/lm5tzkctSwx3AeWCgNt0czA3yIZPE4iwHvLFRXeNEzV9B7cHk4Dd6DvUhqMn63K6VrJon
gtap2b7JTE8ekAtXpR4KMG66fNo5oaFq/oskCo/uRPqbZELN1qpKeMq+dxa5mrGOud2SNAdwoMjt
tWqLlbPAw1KFmGLOYNv2vrBX7TjWhzo69N1AJ2KpcsSLYcvccWy67K2dbzraq/KCkgNBOBKdm6lf
Da5OYj66Zh+dXJHYr/DOstwxgoIqrMgTCvVh6FCqnAZqwbCgFLa972Ju8aVYAcGM155EqIS2Wtuw
ozHpyYTuGDueXiDA01uEbGXNOJZk4fSlxxKXKxD8C+pdBorOawsP4C09sQuzqITPRYmtkMDnfQv6
AKlSprHgYbLv57WfyxZNttOnqWAlFoEJ/EowtVvupmUAy1EYeb7l7wW9qFy4VwPJn2rMYRCZ/YSY
Ku2y1M7MwZWwuWia7V4V2Tgo4T4nDXRIzbs1nbBhrtOqgAd0safTJRionMpxkdfnHYyrNtvicg4n
rQHXfgu9rUJQ9X+U/x+q+HGvGzuFQ9ju3o+rqw6kozqV5UxMcbP3jrSZeZZ+XiwRLI6PxNTT6oMM
a5bteztgJoyDqC+aNJMkasv3eyMw3q9MZ851wRHAt2X0UAPdVsNTf8K7//6fERYcevNhhmjRlCL5
0XzPkDPXXfSbDq4rmnurFnfSqpORzpFpbQPAaxqO+IkNQ5RdLYC+2KekiFYUNIBBNE5nqqKhPNum
7J3wKo2wtYX0P24jLeEW91N4uW/Lrj2mJyoB+TIBtYh4aRhgY+IKCb3VxPLe2BQy9Qn0b5IJ5iVa
zRtmyAOsUXysncmxvzYXDP7KFoFciJolbTCateSmHzHafnN81LDpfW3alC+5y31CzWHKk4a1lARI
SffEksXqemffgUPgiNqi6W5ReOLvESOX3hpVguvaG3ffLAde0w+/pjqTwe17xez8nXwurHD3eKH4
/+nEaOtUOlsDaFZJLieCc706ehTlv+kEzjm879sAoadW//0DnR3xs51Q5+X3xBvI6CZ5o+C01Svo
0nSEAQV332S4xzED1tWLratAIHKPcTmztQ0JLHgZwu4vYEFFMx//GIZSfx+Gzn3NEkHcuLmIDBuC
kHvpuspoZ9ElKuRM79PgKQh+FFclnEpKM9XR/vCC5Y52Gx7q/Ct463G1UNGUw8OsNVhVwYSew6fU
mVvvy19e9Dq8KW0x95dpPnbdr+zy2mF/uxEctuJXS0hW2pLtfTm+cxcoUaRtOC6mz+spr752F+72
1UEGG1TY+3ZCLoYsp6mwu8DiJPNIGIx735gVJleN6fKdAco0vaj1Q9itCBylefzeLk3wIGARXpQr
M3ICPqZsOOQ/wO696zZy0ecfgnBlHqMjP8iMsjbKgVYRVYc7NsH2txpTS+2QhqKAr3jEmgg2+dDL
vyD/RjIP1+jT+LWsfPf+XbKzZz01d/5G2nYwvLvl1uP5PVms14K9cBKty3Wh5NsDuZAVTLOhlp2x
KggRwB/pr6YBJ0L8V5lSIc/DKrXCdmmkHdRyPN71z264xdy4XUSavqXauSMziH1U/D+2pO98Da3J
+Ov0fH2BuIVIVIclmTFPoXgW+fehwZu3ZjoyYQl3RuuKk0jAhq53Td1+2m26K482kP0ozq+E3fgE
G/9DAm9GKHNmb3OQaF6wgdnJqv7FwGMUa6bDZe2v2va4m8BUHV1WmOdYbAmgcc8KHZyQUotOKWac
nM6/LUk8XsLwzTqYKj0B0jblH/7nZ9U+tu5yR1hKqo9rDObxP6STdt02moh810zqggy88GX33l0N
zFUfWjmWfTm2kp5BhivTA79gc/jy7Z3MrvfXVy1Ik9mqUiHsGJ1WgiJxAZwgLlVmzfMBhs5sEsnA
r6TFxuXHNosZOJ5NKmvInKXDDsiC9ZiS9zR3Y+SVxdQDHwsmEy885ZtUzjrNaRQI8h0vA6e7EhM2
1LzNh5Dte56SFrCPbU6yzp9QYx/O4F7ufgPQb67Jc3Pgc0D3Vaq2kCrz3dwcQnfcu3ecYEjfycdD
VT7CSpLy15FgMiWuUH33A2a4YyYsr8xbwRfNayQ7Ymcr0FxbHDp5Xo5zo9F5ZimIN8bYq+eQx7Kj
wuZXREOVTNAf4YVlFYh4UubQesRff7ZLBrmsprQvbFRfq7FqA1NFewOoWIC6FXftOTpK1NUZQXXa
UQYdVDwYmcdtUIa1dnSb+398xD1QzudWotMeagCjWEi4pz1fgMkKQTKFsCzFT1Leesxt+qWVBnS7
lfOXyJPWNjl3jL8U+ZmzoT65qaO1omKkLOTk5XayDvNifWy6pQjwNT8NlyCyjR+V5rcOlcQWclrY
lCu1z9d9PKpCvjhxCuAYjUVgmDEH9RQc+xR0Mhg/nhU144CalXlfvG8ukUMT7arZCqNg3adJidrK
3mkap8UP2GzMS9wF+SwhHzQX30fBOxOvQtMvFjLVScQ2rl4yXeqBIQY+AQ1JCEqFTfQ+AH1BQEtA
yhCWWGQArftTHynzO16LxtS6H8n3fNy9/FAqrvUnt9nULriGd3cyg/Eh5yCr+6686Ago75cjYQ9o
wePzWOP7KYv35rpziOmoRVJeiHZ5VmuxPeBvKAfp+JSP4Qx0IvNwbsD3inVqbgqUUvNzyDCDboTo
Olzr0NT6tz36Gr3DaWlLIbTVOF+0Ia4TcZfWneiyN5hMdOHFPkOWXjDe8RSip8tz2kcmZnHIWh00
QNmLmi/Yj3qn9cu0rZWbml30BIwF2iR25t5ydWKER24El/UrjO6IBgl/mb9RFV9adfZ0F1qxv4zj
Dy7NESnPBkFeDpDyIWq+Qzicl5Te2bWymPbcO7Oc3g92gqAIuwNHXQJAcmSk/N2PtFJ7fqsJtRGV
dz1fsRU0Rsj8DuDvV7GfaYphimO94RXlpb2QpWOuwHKobxuw5VJrhmCWwlvuqjChkNxT40pZQON+
6eZDy3PutXVfqRhvvmrwf4PCk6eO9UE30Xqto9ZeY1Yp2omdSKmEHpOhervVGsU9ThFrBdO9Dg3v
zqJNIcixgaMoUmddRpqIbwqZiZ073xBlh907yQJfU9iqeAX5OlCgjqaibKYzarttB9Y/uhNVA0hp
LiHm/xJukuLmyd/ScuEuKI1mNXNmFIl9OzaclameuvwnKujx6xYckDeOlGU0bZRCsUolSr3P5N1N
+T8LGpzPAOGSU+fVqkLI+l8yuonHB98o9HKGgP0Ey534c9QGepnwfZRp3hmdMKmcDI0SmMDo6Psd
qG/PFxAXt+AtkPHZ8uvv+Da/RWMCKL18GNeR+elJ9ZXIJK6LSAcVqNakotxCTli889ek/FPf1W3u
/ryO7vmYLyHFIgdG9iHO9nSgRnEMi0vyJbX8BW5gmO4EVK4k/S9IB0/fozGsstIN/a60NyuS1E3Y
sph8GwkQjXM7NikGCWbptQzHSCStfD9NIvkt8g03xbxSrYnPNc7qz8SRhRM0HCdnuiClznMHsio1
ueJBSqZrRocbLAG2AFd0TaTtWKwqGecZczWThayQiS77RuTCUH9MhvcQSZ7lQRfG7hdFl35xP4/s
6yhnvfvhG0Iu71H++pqlJSygDNzakr2cXMpXFO5kRiuEat9+76Y0qcSHDFmYdW5C6zbEqCP0aOLs
wKP62Ar/3SRTpOb1b/PIh8qmV0zwFImPov314d/LNaSvq+YT0kgj+zXBRQAvNF4E0g7irGF4rmnH
xh3AneiGqAayk2ClNlUGFVQlnCllIsHzhMJXpOvRlnxNH377zas+u3+QWgU7f/lbdJQkDDMHIvEm
rVIyPyfoy3ZlLvfA+Stk1gQtjv5toKkUx5CNI28nsVyEjaVh4sOAPvq0VGVXDgIaw4dqMzd7B7j8
ofG7W3/u6iLukKLWVLuavzPzD0UG8t9hqxjIBf3sZ0zVZ7UJVS8b+2++/tDbYnuR5cMVG5hCHkcI
hT+IVY0FX1pOGczRDy1wOQ4IhLlYLMoVdKWbDmR/WA2w3+L/skvfjnPc/r0X0wHDVPoDldhgby1t
2CIi2/fvYKlZLpZImE/r/B1O9KND9pU1/4DBxDN/hPjOSG1JBaWiOgV0GVZKwGVnWs9gFuY1QzK7
v2Qg3h/liXT8QoB8/AP2OSbjkr6cCqvMi2bnM5rHpw7NMKK4wmB2pxDtESZrlP5pXVMGz/nD4nMN
DEy0W/MZ298kuaXqb99Qgpba4HIvekDtcw8UJCw25jHw1M80OoVeMpHQqS06KrJNgcVN6TxiBlpn
OTW4ku8JYJ0bsHQmcZ4at8jThnwG1HkMdsOZulW13/Pen8UqPDkm/Gk9lrjOXEHS4F42r1a4gimB
ploilmfzXSUX+bgSliV1JkMVwCcl2YxUQ73rQcfX2CbQdj03S8trNhOL/uWyrakRsDMVIphI0Xvr
PImmPl6lpn+NDhWCBHRP+C+AT8FMdFiD2rlOdq9vyuTr8tjDklOkg7IT26yUsVCgnWYXWTZEGNNq
Zdp9jp+NNUHnKaUkpAtFCD/bab4cBVN9tzKAE+jJH3c/78UxcJo2tuEGG6yFeDzTi+5Aj2GU3UFj
BQVigJYVd2TvwnGl3/mCev3iofqb8sOphN2Fl97W/S1LNGgmLBL0XWd+YZ9hONq1JLNE7VI6+x/6
dfEo0WyQC2UhCzYeVmvALCiREpTpmX/+gP8Xq+E4/Q79YJPnbIM7w07h6O5OAzyJAM0Fup/HjvwN
l1M7Sm8MNAtFqgu/5j8Sof3oxWgBXeic/XAb2zEbWeWZpdWm8NeHoda8DkNx7sfnN3D0zO62V2rU
RdW01irg+CP21wK3JM2VDzIIjT+0i70Ir/K0Rxzo7y/wi1WlzTNzoHOJr5BkeJTxA/1QDj8cgjo+
wDXM1luw5RSQiS7yATf/zZ2ludjwHUT4OF5fGTlzhDRLfLf9Oin8JYdkAziKNR+5MXuzdwnuQjJF
UX4dne9HXu+gRPoZlE3JoRs+XpxZC5ekiioJAHw/nav3ge8Pr8ij7LaQDVgQ+uLVi2NPfkNkxTSs
hoRae7zcB86TIxHQBYOf4hgNFnCdp7Sj8b0AxV0cQVBJeRTuZ0QXHw2/46WZhzm9kzRyJ4IT0DUY
7Ora8BkNUVS+tXUegARYEHx5krxjSC8kLUHYqAxmcmR6yemLShjW1UMiCDLi4aVidC6ciVaFqW/T
oqw3bJuDkv5WsLatEsejdLa7AELvJIrNO4+nfi4swkAypw5VBq+C16a4Ueup3zZ8LlYk93LUBUI6
wToURY6t6ALS8CXHZTD76GQ028Mgy5e6zeUqnf5KyjVyrtFSP5yzCgOPhtjl/AOAgDmEZs7MRheP
BP827IpSzWkPI0cC+A0NYWoSgtv/X9ihRXmECi954FGckzu0LjY7hccTfQcsJtQBJ0iAhSkcx8I0
H+ZHetlzsVTJx0TRZ0kHbywt+cG0SmgingzhCOIx1/2H4UrOz7JOkLBeNWNCayOwkFqcLxraP1y9
sbuF/wJ9p65XTwboEHsqm3wBq9qAyiN+2WSq8P1Qdb3NPY+BnpjHDHERoYogos8F9AzKoyc34j6K
Hiu72Z8+xQoodcncyST6xoXkieZQ+GbdAFewSA957x7fO7eGRgUQ4o0dmXEW1U0xBpeFkrYjw01V
m/V0WVZQta0LfK82hwe/Yyi7TkVu4HET4pSy82QiE7Y3K87JeDNosshWYFHiv3wH7Abah8c/Kec9
H3bwWaw6vRwu1nP3H04WKWTKhLZuZg12adWtDNWSUzLRYRwoo/QAPLGoa4mOo4cOXfABtKBAX8Tr
YOTda9VGUcXMKgMkmbMSnLW5/2HKWjHnJf42Fwc4vhGxLogGoKW7qenK65OesEoNG3lTzKOjZGQj
BGEh4qKg4ulE/NbWT5bLuFmBNp0LG9PX4DfjnUZUUcpibGXwtyp8PQS9QNEXAfocsmPc3eY2+LZn
uqkhlLoupbDBIrSrQeN/8/vUGxcr64plD+m4SD7yhmq/oCrL5vvoK1+nohw0MYmhPyyVtOoqR2xz
9rrTZfyvbcZvsHI2IiC1pzH20Lw082qK8L50hF3roXYN9CXia/9QG128UH4+JlqJ6qcFzewoOcVO
RtZ63iygsxbGbo8hzm7V7Eg4UGQ+Zm+mOyJW2Bq0CGVXabmoMWyn6kuSDHwKwPxaRgoZuySkgFVb
cn4ozo7AaD09J0BqiKTOtXX5nUpQtgvLW8JvoeHAturRIH673RTvpe6UDHca36DV8rc72c5e0a23
oY4AtpzCjMyWnuaTnM+GwuH2T8P0uLqklPGgnLwcQ/2PCSc5+x/h3go+tlNXLAQN7dNkdY8nHkf7
eSOxzd2f63KSeIIrCqwHyL1/ZME7S1LmBTZiQtK5YzcwUTARtEz9K1RU6vKWyXh2PSnPGPC/nRhX
oN5m8t+XgQelTjRHS2XY/9lNErYufU3lfA9JQU7oumKnoLrB9Vygq7ARd7pZq4ho7ycTGy7SjLoq
AKRXubYGfqQ7biOhWn1GyXFqw+3w2xJ8B/mIOnIv7OCTS8SixCmlCAhi67FVZvBMnhlgPVO16eVe
9o/NvhOEY7QUO8QCvJ5Rks1dWjGWbSOKn5v2dS5yBf3stY1PrcHjbtDynn0Fv0ejk2N3TfKr3oXt
yYR2XrbiXUa12cCuPTKk9DJEGavWi4ofZe79r0ye7hP2exRXxMjbH6kmErRgBTL+ETw4zo83hhNU
k0IhYH+bjQKNl1Nl6voPT/QOP8xhcene2V2FoCcfApg+8yBbDi3Lb0CyEby8XGC7DbP6lgzz/2DC
ntG48V57SHNqmjxKwS88tuggYp4zy5/ZQ60JXSAEE/M5xHZSkSA7TRgfD839lg6n/h7WjSHqo8f8
fVdxnnQY/8rM7LxY2L0lHVtWFCVjMrgv+vhXdZzs9wkfdTpGH8JbdOCo13l0M9n7aZUsvbggOip5
YTIIa9Xx28ngthI0nxGcGwg/9BYsHc7nojodwNC7IF8i+wBtZYVKAGQmYDn15Ka/a9nsnhhfsFaI
9gbhrpD40Ga5lz3p/gTo3BXXDgE5fc4R6aVCy2dbX/hS9sMUnOmbg7i3YRNwpIRcKxYLj+vPgYJo
KxTupgVlyj4yy76WRSW6rm3iVGfgtUYPe5qkG+TKNiDgVUNYoe4tVeN1OFg7tBaDg3PIHn5hRWHI
BChMYdca2SrLlmnRkOJExtKR9SOHyqGG/SQ6oti3kE2V6DKp/4sx0/Gtzi/2FJmCheENvXUDEizB
M9caGyWY0p3Aa+d1y3d3xRc2/REF8VcCECKTGxcp/u4n2c/PhfFt4XDOhyOayPZK+FJb/kg2yOKk
QwLH9Ys7RoPhXSgbHsV4oKGI7SiGss6YO58rQeKj8Pcm3T0Zf8gYaq31JCOjp1hH+BGcpm/Z/9le
ph3O0RHFNX2LGBAXMsKibwc85Yb/PPqxn6O73WXN8fP5QiNizbNCNTkDTrw15OJADXgx1kUlmaSy
nrJFEbFms8X2OPzISiwXdCYX2nYIu/d1DXsu4pH8ysGTAaHV/YajspQlaDMgtSxjx6iZikJISIS7
JMaIZvFSE8whiKYZ6NP0YWpHOl/LV6/aO7TxJADe5knd67vHVehHrdrOY5Pb9fBnvAtRmPJ1SyFm
bqtKLm1ghzku7AVzWoW/uivZNesHkaOUdvlEEjiWz3iElRgW767u3jnTyhw8xx4djzyyLOxelZ6L
N8r/aAc7d47CrADx3OKNLl80PbhrkoNoeDdFe7cWbeZ0a6IEoIy0MJ9faKU3QhvZis+iP2XZUwre
OAaG50J/FkwteO1/a1WMe5YhERfCS7SGjutDqKBFWRESIZkhPr9xJGfvhWe1VlpobVeEVabVmqwn
yD/h6cjKGCJpLdVo3FTBXXQ7fALiCuC2WgqRSqPEFRfAmTALasSiJhx6Aywp07MkvOGp5zSfxFK0
Zz6Yeooqp93Q6jQ/kaOe6fs+x3Icimla3sq8pEu9TA06NjzgNVA+Y8IfAIZ8JyumWePUhkoy8ozQ
JcNH8dcekb00oARefiWk+mhCOJztHAT4my1BQF03xJ1trmIGWZ3oolbDt58jMvxuvwBgKGIFkCi5
a2YlelCzIlpcvB+VpF08Pc5WFCyaen5yjFRmQSX411tcNJ5pnTV7rChCIHNy5K7f7qqA+Y3ab3Bc
BDU85KsTCUXNSGwgDy3qsddG7h9vNtzORB7GstHFa280cp2TnTI+K5eFJR3w8bJ02xBRVK0r3YoX
6M5QyHNR3xfIBPqXQ5P6zx4TN56tNifw//vU6GUut8MoGU85N8yW/C0J8/ZDhIjgMPDWQz76uSdC
IzPrsXsEfMTwIt9FEeILNCFgC/wtwJTxRR4sLGXp/tM4I1PtsIIbO9I81kgbHsdgvvnaGZwSTfKx
3fTT+CDVyNgboC/6mSikl3QJQN89tFE0xP+fABFaC8agAUsmNChF1lIdiKB9/pKLnyGc+UcudSTA
NGm5++shUHzUnHtyHL1oXIJl8wYc+tJTJgvbMlbM7Iqh9LLVE/lRf34hMzxuyaPz623u1yKKAibQ
4vQ2HF7YMUSXjdxxobbPF5yQLJo+Z5K+6+dDWZ6M2W6p1BCJ0hwyAJtKvMK8sXmoQ0lI6M5jOk9g
32Pk514Mvxa0T038t/lGabPCNjb7/HMo/Sa1H2kbBdlcRqr/T4e5iN8v+/zN55aPyakinJXY3lnB
53FoAQot+LeBkM5CAZVfsdNrcAJOA8bPG23c9swHYzNcTD0S+jRHhRfgBMr9L/zoOQ2xPXHVSiad
NcbAhKYBKoTopuXiWqP/3Eaus9fveRwidChLEleapw0DSYbrvWwBjpy7fu/SoQdyFWj25CyhLS3G
DlkU+Sqt83iEliM+CZ9dB1IbkaBXl7q+temXe7Ss6X3t0TQS4GTs36rQ8aGf7rOcp03q+YQY2QoO
pjqp2QUBcdvhfZXo0Gq1N6m4MafCWFR6fqiUp6bvT3KnWbkdj2fdswsgkopy0BGWQGMUPhBO1F7y
bdg9DkpOd4ugpiO5d70999hwOuffLzqs7uSalJB7VE6du26NVIZ1XN0wpOCbZqUdPp1SVcLtZY43
RjhuRtCMAO8iRjNv9bK2Vy2l9yjAWqboFWiJoBNYA1lwSSw539d/4p//fOvtnKsqnaPMp76X4MZf
2zgYhpl+rB59o87EsMKze1HE+TtxpWP5D0rSE6f4lGTLYcXHFHZOyCKegklC0bzuwOaS6EZCZTi+
HMXkCIT2ObKbdfoKusfzh+tCocK47MLRedDLH0dHKtg0N+qR3qBDjUTmDP6r2lnO10pGg+WfFFJJ
K1rk4jvmf7QCphXR309+ItzpYxJbJ4VlxPuGZHjMSwWovGnRTpA5s0e1+1rpzghMyImykHIbM5Ht
gkIoko1KkRRk9qn7Pjzhzoxr93KRAGDi2SaUHLq/ar/k0M823zxvhzGL3H+7uAu5GdSinHqupo+q
gsU30rOMUKlnWcqaa9nsyNCERYh635k7WpaJkzUrQBwBocP1/qGN39jUd+ncwE9rQcy0iLy6/qf/
9ToQb3f3obtSlkOqpmzus6sU/wewwewBXAP/I+DqkmyhJMcC2THiMrypQCx6CfcLJ08Umr+ov3GJ
oDgJWGJiumkPNE/ctJNvlS52sXmd9mvy4WS3VVpIIoA+Rc9x/T0o6+PitBN6fn8l9TB4zignChXP
UevtdQ/0BWUvEa6/GQtqdGtUBi4sXdK7Hvrnfgpzao2gwWwWcu1WgyXBBEJX7OxCLMUTLr9Ho64n
linIpmyZll5T4TPBkuS7k2wq4yVjmslJMLvpCdy9HEHSL5Ae1IZye4uMrJfYxHr9qRTk9r0PqH6D
wym8ly3Zlept7alMWkeGAyOJJtLQBH+lD4Gh998+Gyyb8rLW96xBWN2nS17yJ6zckk+bsaH9YfY8
U7Pi/F2xEcdD6p2SO7UJjfRo52bXVhxEJsngDJYU+NUAbk2aOAQS47aDpw1oXLUgFbuBuGqK1J8W
xZP9rJAELohUUqVXrL00peGGtMYqvRjjdHWq9VdU3fdr7Ssm7+vx+edRjGZ9OuY4kZs18iJ31Fzb
+DuDBq1f5gIvfzGYb1aByJr3O1ViPd8Ndqj+kL0CdTY91sFcbjgzBI9gVDajt/7Nf7NU7B0yeXPK
KePKYH5462H5Kscy+MeBe5Z/nCOaa0O/PakXas+jxajKm19e5kEDJl7OJZtH4brKb3eu7B3CIEXw
HBcJRkpG+QffhX0qtFzzP+ClJvjnKs4oA5TX0+Gtszqkp8qK3XnQNuEsVsaHrcWQEf/V7MUV5e5B
mr34orkbloP9BuCpYyBgrx5cJpwFS0RqniubedHTaTJmEfxC5D7B5gVzn/4Dr6BVRAqgiEwgMCv7
JjziRdhVL37Wrj3XJkTxaogO5AVaoJ1rcIN5rUTC+mDd6SvX2nLuJOwPRfTveHwQrQgRLkTFS9JA
KyFzwOxsqdAGU+Y23yazCdU7AsP0IG+cErrZF9+5o95IgSXpb7+KYc+vWK/yRSmXFbEj6OSZpVLY
EZeXFfs2cOMDJEr4KYoqjmioqTuSJ2j06UBe1XDbI0ctg8KL6DTg9XGwa+n3zi4Ylo0k26s6oVDx
MIdSWsrvkX3a7HYWKmVbbqkIkO4QGll/JHwJaTuWmRul8IFkONJOusit7R75gKCGscoC9CDvLyfk
j7EvVLO3BxYWpufGzKnFmHNn35H1Y1ewwgzK7Gu9hDaJL+Ey8sd312eNQ606IJP3rUmDEprF59sj
d8TzwccMc0DrGxdElgDx2D8WvjyTsZjcITigjmyayyQVJR6/OE32Ky/snvmKEsxCHGvVG27Lz3ec
XfUtMzyc1y4WBnDdphcY3sAnea6Dx6QzGLTje+3xxhnF2t3M6vlVrzSYlXv72dJ/0FJrM9m1lPON
6NXfjnj0FA8PG+nuRS3FfkzyT93TzOXYNLB9bydmRsxom1xhNlAeDAalRGlqyaI2C6VH2/ML5D4X
YBVuRVFUD/VLuk5BpgUEFWjRqxAVx4clRLsQhbr9QTdxljPRYbT4tXrSHFC+pFJDY6MMIGrMM1N8
Vb/YRHLrJW7NWPQDHKySApM0rlJIjem5xJqRCjxRp2VLpEEhYt5y2mrZ8ZWCoK26uHyHTgQWTr5m
vjxq8RxaEFHnL8Ys21YPpDMl+DJM9fetjuk85pzfP3W8v7vLO16k615sOpwjTMEsGPs4Et4fsvwn
oJJ5Mwxnq4LYJ84bbcooo6XRfollKHczBEZwch/x3znUXTSJF10ecsBwqQY4fpc1eGzj9gLevzIU
uBOnhX4ttgAcLiY0UQQNqXJr9nh4tByjEc99bRB5ujyE4Te/B8F26PDgr6SJ6yyHQish6qUDTnwh
78KBkRT1P7wWh1mUwrhzjgxoiCV7vUKPbNtFjFc7uM2evFsLnHzFVI7tLjAOG7ym6uyw2hJqr9hf
kRlG6oFwZKuE+j7q8VjN7lvqxSrYhVud3P025UfCt8zouFUzdNUPT+3h9zRq28d6ThOLB09h7rvO
+JD9gRFzSSWZHGXyaogNS9QJ6wxTYqtbg1ogBDSHEZrPHSFeC6zV3y0NSrMNMpDeG65Lh9gYBwws
FCaWiWDqn7fqnZR//0mg+Se7sMG4pyB0tmz1WZ+uIisHqrySOeZ9uriH8mbnY9P5HHYm3oLmnt46
Pm8KW+dQwS95sK4AAP5AJlJdLlV32n7IKyyOkhJ7trN38hwRdN40b8mjPttp2g3ABHOvn9OYiA3u
vEQgl3A3Y1cVj2NIj745XNHSDPmeQXZL0V5uHI2OA2BKfBDcT3CxP6mPoDut2VLdW/6lta3wFVYt
bUff/AzTfNKlmgaqc5DrqQajRPbZB1nG5uu+032SSc6Np3O4brnv66EogZT12iJqTC/3i4YOH37I
DzwjSxlV9tBWAMFjGUTzoMl1d9Zim3T7FhIJAtrsPEnI8OD229Vq2zIUY0tK9SC0sJ5R/utors1l
vrPlOqG1vxD+ix27O8SAOtPGLTyrVNp5TfITmosNkgr+xuOw/5ZBjNBqerrZgaE96qGb421umnL2
iSHlMsZQRg6hRmsMB/T7x2rGpWsOgo7uiGVDoqAiEY5SYxFwJkmRmF93TgJnMXhoAVPlwMH/Id2A
ZgXVb2+LVsybDZtFjcMW7Yxy2XBzD0PWnKbhpmGZdNKOQ3SWselUgKmuTpI6/E9s8iHpQPG8hhAM
G9czg9/PlbMfdznaCA3QdHnzc3WxUaN88DsrahYc8QrXSHGSu5w0IFVeBAzh20cbxfrRP9iyoxre
SxX0dXC4iiGU14cKfyCoFgxTbnSgQ1S8t4TbGAtt7ZtMdpl40Y2R78Cwib774MHxagpItvSoZaqp
QzHqHt/itBtb21PJvTDTId9Im6dGqfOlo83orNGhkRVPTOQehgyRmUTmTGzDeYCQexxoz6TjFGQZ
quZszry030IdRcM4E+UYq1eIbsIzgcgZbm0tnSjQ8++3E4LrFsaWJqqArsULDyhL6ILWfLQVx93g
qH9NSRAY+aT6dPPNJzU+TauogSGYF8Eum5u5rxSZ6Xp25sSVsYETb3mug4r4SNVWx2zFPicMST+A
5BIE6TddAF/nJ/JCKTQ231Y4WVIWZ0Wgt+SCPTjX3oy6i+EJj4ZoBnwhqNbKF5tATLexL2OgeSWg
KY5f5Nh38BH0mA8qvCxB4sYzl2CslBIQOKeUfiqjRSycVcUmD2foZuGXdKA7sEyOxmxekRne/P/u
1+9xEhxhNHROE2DMKC3thpOsyT+jHeQK6fanyTWqV3RUWSSsCHMqj+3dOR8rKd8Wdg30m9ZgBVQ7
I4VuZ/7P3BGJVTC9vZpL/tuHYnxvsuowcYSd8Q2BK0RsXF2PF2YvfHH10YAt76e6kJZ6xLJ31Nfk
QVo971k6+/3RlLK66v3ZzuGGvSTzAepNcTfA4XoL28gPL2Xvexb/75ypHxFKoYuWoXRy0W5gvUKG
xjJSEzIDggEsS9QbBvZolH7KTJxFdqLwZ3cL/sZb4S/eQ6mJsX8GMq9YhsNX4+9HkmTBWRsupIlm
6EeQYxxTGlxw6r+Yge8RwVPG6LOS4+2ZROI4znY74JhHu0A7aX+mHU2HZfCyZuX78R76+P9/TxOV
G7aa+bUuTl+oOKchOKaWhWsm0ptk7za1bIfLFtoPONX7Hyfk6M/Uj17Wwx5qbKkuv9XzQP/poIlo
Rlc6AetAmKsATygt9sUIhUvacP1NRzxdQalIHvg9+nxI2j8CecjS+V+IAdsQWm3nNGwJBlxN0J8F
TIePDbu4NgmIQp/K55gr5PW4B4K6CNQr7Xh91xCg5BF9RbpEpVXzJ7gyp3oGzfbIZpJt0DEgCPiL
lNXhXjZouhCVSl71B0VuDDZU1R6LHKezswu6Q3y3AoQMBesY9HvDThTRIxm8W52icPi0p30Nc7Yx
Pg8rGbIYRYusS5rMH4T1/qrW7yXltihj8aVk/tlNRXq1V/wooe7k9Anrkbsnth17ybcmzTlI9tXy
km28FzwCr6uBpKvMVr7hrUjPRH5FLvmla9izbvR5FNCCQiZILeddL6qtfpp+6y4RQdkFSgbZt/Jn
tl44y0tIAk6FUbZzK36AqkZ3HuYji1OgOlNetaXFI6ipA42ubN3rAzUD2l3LhnP/Map1twR54vt5
IXAejYW56wt46NBpRo3RrvU22e0oCtwwZLBUZljkwb3GCH0/uLksUnTbJTk8/eAGFjB2OjGk8KSI
AuXsJx+lg39DkeCpgPshR9pVDW6ZPIKzZNKSDOz9gS+XnRyCnJhbeLMHMhmF+fo316SZfEjgSgnQ
F3xzYdCDo9MaWyVMGU9123V5zBYXMpbdUuJ0zcXmYZj1MQ+6BkjENFV0mbvsnR3CBI9XSWIW4ioc
+Ku6SYZudB3NQgYl7+jglKiyBQu0w9uOAzDOzD8F/Ht85XMKsOJx8UQUQfIXSrpJHxW6UtRpfRET
MFGVON7x415fJ+jeOT6H9rbDSfEtRfSlByrvYPrN9sbk/OlnorQckUSmbpeErTeFLXAQIPOEo+qZ
/ILuxVXElHSmfPZlyN/hP0Of/u9UG9OXS2Uf8EHNTvykHYOzBQbsdoKC2tYmeliv8LKTWy0UJ23Y
AkiA277vmwum7mjFBLIpxl9+7orKfhDZu1Cmn9HIUZXz/ZYbcXeRh4BSzSnGBt9RK65haCxAyeT6
hfiTKXuH+ojdDjfTpCjcnld2A/Uuc209nVQw7E4xGZ8qyQ5+I8Z/60+XvcNRWfApdTtk8y7Byhug
mG8f7+3mOTHDVtewikVhW5W49LcUu1Wj2vnrmwmUyd6lrgiZgeEW4XMm8fdyS/Mvm8SzAf5ywDwt
0gnxh0ObGWeSXTGmKQKhzc9AcYmaa6AFXVtOjDP0glZOCH4lk7a+6MwiK4DHUjHX9gCUKcvJiARe
WBTrAbCe06J5oGbR2lUfuoGJYMRsZr5mhoAA5OgKKNS6A2dCpZUNcdqlpsz14uycexqSyKtB2xsv
0CN6GHw1r7Gcroh2RKE0QMy9Y6D/icbRCo2wgKCDp/yTy7Cs0N8B0mvpgnrp/m67yEoq6m+RMgOy
m3v4hiEsoOFNesa3ZfKiuIA90wpHNJoq7TOeJtymQ4o3+UzdZw2nrT5B8JnExyiVR9VBdVArFH6K
ZbNAJkJMJUGbQGvCt7g3MAI3Jw2zkSM5W6hJGFXJaEteIkVwYXFinj9ekwtoU2cF8QprsdcJZiiF
ckWUvOE7EeUYjEYaQQ6ySqevYDvBxSBrEXGLIG8T+A3/FtzjMTKvhVeuJKMV4CigEo4nZy9r8Xmk
SETDTJabGE5oIRWcUxr/JQ96Hz0F1kTbYwa+TXNqGrt0c59jnIGXAjJmenxJW3jBP5wLO4MzR+P9
vxpvy5onKYnuP42tOlTY4w2bxm/tPE/EE7f2rKihW7ZD8LmuXDoFBE8P7xjOQBX2941sC7MkYuKE
/0Pn0ro89cAIwjJJ32NA9f/RrU/vUV9Xqk/INKOUalgk1jYiDgQs/JOpsdS4yhfT/bAerFmXxbrP
omr4Wcc/HY01QzyNJnufv99hLOIDbJ31VKOBbwT0DB1kMHvWf3qDSJSkxMgZDTogL8/ZbcO21n4y
AQlbCpzaJipWArQsbSNeDhBtTikGx38wr/4BNX/EHn7rQ7FWZdC0u8dpciMKFTUImNEYtAD2A1W0
EoSOfLg7ihXpVZe7TZ0MOqHwfUskLkZY/35fYV5Z2zkw+UOdz5iEVF5yhjGdGTja8s2csV7VhP5M
qf/ajqNsalR/UnT8lcTPU7rRRHhRCDSsDE1xpGj3lSZdS1ZY7zdSbtK5AccB7fE6KSi0VZnjUvtx
CKwp8ewKIGe90Go07H4KcJeVHdMSwFiTKI++sNkkZfN6eTiGpvFWPVQfK7/+rCsWYCi8LDMFBKLO
Q1hV8/gX6eoc0hVBoTahbpP5wbiEmjMeh8sWrrglAPJ3bsJ/mn/ZSAKcnPoxrkwyWLxZPn60pcYU
rpVDRZZD/QxkNCxxqmtddVuEEyXmpT8mVRXok55Xn6uxgkNlZ3TlnHFhSkXcAA74ny0diTjd2efK
5qgnvXIDnOIVIODftXG9RJOLrqJUlNY+XI0qxMtNVN886BvqyiomOt/PNg1Y8X2BQXGFJC6lu9HU
7zWnT428lsd/sRg4RZDEggyvXU4whM26NDdJL/P1UQk/KbQd7QqJmk2vlg1ZvlyYYgscg6956Esf
uJilB19e5QpwkUcOsjjppYVW+0yIXkJ77crKvBmY4caRHDYBBJmbu1dkEw6LxDTjTGBOE+9f96gr
8OAWiuxnMW8gKcsNKux6dJcdCJPPus8Ie+uMQ6qmkQedJxJdcCbYDB1iyrzNlujddhKbW8G5O+UQ
omTJilTTMnxeXHagqPiqcq5NYUAGuWouYw9DmoXcyZ7Abe0SutxFNbwuxcR2JjOUZpYie8gwlQm3
LHMjgNeFOcxXNlAyorCrerZaLJsNeiOQ4E7gc9tzUpSjXVc27qkJlV/jIDYPJutnp7hJsNrO+S2d
M8ndXThuvGsCgGhSWfc1wUk/JDQUeHXevATPEEY1vR++n4IVLKDNtGlRPhz0KZc96ihpDG3GWc72
/Qh+3W+XwqXqWRETHHdI7uTc5fW9ARZPOlB+n7SaDl7QObgTr+N1x9uFuXR020Ro55H56u6yKJ9z
gMFYbNNAvyfQ2QVhYwrdQgy+BcS5EKMZ38L0Ct43hy9BP5BDHCthHIyZHccFNOZhiFewqClKpLAM
YZaHG4c6XFkZW1tra8IBOvwMchI3179eMj7FcsWzA8wDb853PLDaM/Cf9JHSs/Gv6mwXo0BHzn5u
HBFAWB2/h3ng6XTrqNvfs7AX3KD4/169uZUdsv1tSLVQk6XdnFmocMM5RwKQTw1Fz7Tirr8EbkfN
k6e3vUISLyorJB95vvs83m5aU4aYbmBNEXK+Q1AuQZhPFbL7k1dzHC5KVX+Y98ggB7slanfgbbk3
frEX6sJcR5PcwzbiVaJfnyL6BCAKeyHjH/AVKVHUi0OZnp4isfb2Vzm1lUwg1D9HDIZ4pt3hN1zG
KZu7S56os0H8D6uGWDT2LozWFPc+yE/KQdTOHsk3RjJKQ745RIoi1DrBwmVHAq6oD5FUE+Fxoq3k
vaxILYMGgkH6KA+Thsd1EKzwryJc/tVRN+wumQGKTpCqM08V0JXusEmBAO7cKTWdDDvAqTnUt1ew
jVdVfdI4xeJuwv062rzwthAF7YlY92dazlkZhAieOVd0tdVca9SnU//Kthr9f0pYEC6KeaIriCNk
lM9rGQccSh2gQ1x0pYzRSrn8h39B26fXBdTbYQ6vGluzTLKSCSfmg1V/5XbwQ+Edp+Sx8NIgXeU8
B4FsHXTjO3ehXMzDfNDiJNB9Lap1FsDLrxK6VP2snZQHFZMpXRwXIxn14ryuNELZ6TV1KzugTfKk
3WzRovFa+OE3Okd0Y2WQiQtr9tsLA2+n7YUyITl/93Szd4krAolsezKHBaFWvLrTBD4JfVSRi34L
BLxe+vkMvf0xLQWJd3DjuvZh/2o1tlqz/JFB4RUCluZD84qUbpsVTVIcE5jkR3VNx7P6H2D5yuF9
tU1S42Fi0Bm/nWrGRFJYpOuO010I+lIp7oTgu0hb15U7qM5HjqcYlUd73DlJ4Zpt1tihxSYPvnVo
dAKQ9pSpcJZupbwAIF262gyaIQAeoM7VaoD3jkzCKGzuezAOnvDI9DGGM29h4ouFx/xWK2wvR0+T
EAf1p1Hxgfn7PtA4HMBm8LwjBnW7Dgrzx1P5Lv31qEViaE5xT90CL6nZXwb5Dv/D1ukAaWQIir+h
A39Sf2si+h6YIieY3XTz4IgnAcpLwVzSxFsHQnqYclH8SDmZ9gX/j8yMqsodak2ZsqynCaff/Vap
sGaj4uE9VCPQTOQIoVczd4gHGwdLIw+KsBD7qnvFyD34LPcf6bAFVABZgCE7mtsnu03jjDQqGiPM
MAimLsHfZT8ewKPjvhgsLDKU/2lAcwWF/KXo8KDfNgcR3OpPNt53ccLQ8zG5o3VZ3FqlrjMwfn38
jVNFa6keV4yd/Cebrrmp3uxklkJdD1MPbOm2Dprfc1JNFueWnUFo5ktIVakzCT2IRf3Udqa2HXH/
Cg/RkazWr2cMdX24Op3LU9ikNbFKbdYor1BIZYI7flxjPyvFH1dcXidbRI0XIZzET1ESvNo7F4s3
HHYKc0Gz5gdVtUBZhzwWq0QKi/K/U79rMmUUlu6UBTD6asHOeovd3CTbjm7FXn6zl9PyQW08YbIL
RoCw15xw7COBryTVrrjK9h9WGExokSxot7drJTvbWgvbIFkZQr7AgSrImJHTkAzSbaqnsO3XGYyM
edxeu9wh/zg/dGUs3QBHXoyeHR1rp0LacZFM6SSrRZmJI5HZKzjS+VvMX4wiFzaWhjt9p3Es5IfY
ciJW+dz5WxkuGLmBv//eC21jMKjvW4MaviJHbRbkT3Gd1ZGAw56cXYfjRMlLTPfbWibhAjPCVk8h
SXgEBc1elM/PzvpnSAmjMYkqUkH6bTHlOIyBb4cn2KeWElMxtep0rqkdz+5ugFUTXAGGHPxgaEC1
cJISZvhmrzoSgwsGe8O2XJwX2xBlmrCCsl5xCWtnp6tE+WgHZfddK4AyJNbvSaSd1unJ0KCce3jl
ldkgt/O/ZUE1TmOmhdnK6qG0Cxt03n9Bn9flqgWABg4i4sKZ5JW4uOiBT0tSdV8l4Ny6sKfciyI1
ec9Mpktqly962yNMsCbmA2CUM/F5Q/TUB63oDLfwwpkeCQzGqXOKNi5eZso6kwKC634DnfL3M8bI
cZeBNqbDB4gTXaQh1RSzicLvVx2+daVvsHRToYxAfu5KtwB50/BZgCV61VmMLInEEYk/aVtWEszc
iLicBAusEsLco6El6qZFkTHxIHTnhI9txr6BF0Fwy38/nJlR3+r+q/mFIRTN5nO5CMb904GhgIgK
dN5xPChsxQedKEj8jRnVT0Y/LLxvzjKQ00AoMHlSQHLYLIfBNEv5lEkvCydqk59cFOa7ltOFZiSa
pZtHCs+9nTfiXl51bkcfWoM0whMR8IoJdYN8P+9zPU5PBVLeDH6iXek4ouFCyN9jq8nuhsh1swWk
N4hzd1jv5dLhvnpVizOBNxM2rcPv9aZvJGZib9MpzwxY6fNliKrmStlnpllVpPFUyy8in31LPv31
nsJz3pR3+JVCkJ/ghWe6S7q2/tnesIW0ysI+QqmrzKWoXMchyYzURr49AFx1SN5cyI+JUM2IFZnW
feSkjAsmP86C+fvRrwu+ede1lMFOnZHEfCW65qrPzqERtgEPoJqfQ5u+YNQFO+Ir6oCRQiP6MlxR
UpuyRntDVKHVn9m7NQINEzFmUW6nnBJlHU8vQlJO7s7ErzjsrbK5yPlahP5VZiYdfBwlzQ/28csY
ogf5oQS83Rec6FCTT87Ktl2VwTGKgAmkgFRO4pYpUm4JPkjfENqO851QjfgkPLZ5SMwuAw6tp2un
k0wvgPMxpUZ2uZn9mD8bZPJNrN78FDeboHPNrGBq3o1V7+wJK1aiYZeMU8m5gYvfaP3IGu4UV+uK
wil7vCEjaDchEZgcojDgXLEDB5LrAzCNzbwTg91SyLMclhW/C60pULGIeY1m+wm1XRKOTwxUkL81
mZ0CyburPPy532HQSMA2rp5XEphho1lhq+AizNJp9aXNQSMoAbgGoKS+kS6E3TL50zRtGG3eMNkx
61Pech5ws1SCfYGdMRUbRa+gT9Uja51LvObq2ZXERAzIPPZNI56OowciuRni4H3BVPMog4mssM9t
Yi+VYyytAGcq9DokJciiIQpDq6P5EkqlTpz2KxN81p1hkiq1nNrkZ1igizLFq1lJheu9AP3tHyDB
NJMC3xGaK/mJsH4Y5Oji9rYtrf0Fy2Lgu+jv0oig4nVmifKL4kqR61JW7P5tRxjVSbl1Vi76kshL
0uH+3K+/jRyZz4gayqTOyI8jh4C2a2Mzz4kK2+QnNd9/MrbN8wlVNyxbYp6XclFgBVKTgvw8UYy9
eO9G085t8xo7gGTdu+HIBbspuboJ2kQNUFNSQqH+OXvHwqArfWTCU0j8cGcljIIKznctW5YgEBmi
YL5MOBNb9VuIKErlrH3LH082mcJOTdGjcm8dxRSEvQQsU2WGVdQ3+6830pDZQ9qZVGfMGXq/EycS
YMncUr1rmQE9noZ14ESfAN0Hv2uXoS/C7UKOcmXSQVbiI8nRTeyKI8O5svFd9eNF0gzK75MNaRPH
/Fi3uMAYVFSdyjYedIGj58dWCUVKcfgf0y89wpi3dq61iBiy8LHyo6gJAhlBKe7Gq0VzjfBGxBRm
JzLl/s6wnXCfY+tMc7adE8BDXFSfHmUSzx1PqbgqHMwx31N0Txd3v1VYAZb+PJASqdR4NwOLlk57
lYj1BVUijGyeHPWxBEN4iDlwRjE7s+TXrOLUTx8gDNZpFXpMZ87e76t0xykSWmjGeZSUrXYJ8Vy6
4MOZQkrcbZSdf+6YSw8R/xgKdYFEHAkBKcKCSLeRHaZVxMgRnTfYJWdrD0GBAM2A3b5ud0LzRZyR
aHSZoX9j7FSGW/6bpbdy306z344M+stfhjuG81AaLFqD6pQyGTOBWb2V0drdIM0ogecUo/2XNxDr
KcMGvkPN7BtlJ8dj5l9MoqJR+lVhqMetG5CtRWwri7lH9CvYuwOOimY0MZF3YdXQJdbVJFxg9zzO
NqgOwNyDRuGNaf+AJapYnLSgekxsKAA9jtdejFccB0Sy4zPRvUeWr34kXvnPzXOj4N1ptacHN6Q8
HnfHOdfrhjoQ82pgZJ+v9F9fMnkXNEAJOiJJJZQ7xyjcnWoqoRLeU1VinfeDYu7zI4QUc5uYMq35
YKhKdK8f0UdEIF64dVEyJQKDRV6iyNut0/5SkKfDu+Vnc0z9aWSdeiYBo0op+2cs3uGPIXh2vIOU
3HzMX2UQRDXifkh30q0ggWWUgDCroZME2Q8FRASEjXJq//hMrMX9UmBmzKjo5IoeQsKxZzcA2t3h
mt6ZfIddC94h6PnHwQCPTvcNjugvEMCzXu3stXK5X2xlJIltEpDcJ2BhMiz5ivE6Mrz2NIkXlxM2
NC7cGASM2ejenhOXouVoDAYWhaY5CTcxUT27Gjtx+zetlxt15gC9uuyixJMBjz6M1jjul9htqRnq
GOzuitatgFey/SVKkJDYXpZbAqoMEn+ObrcvFRvtLfhyas4FNbL+ugNJZH29ykI/GyA2All5TeUS
jLV91ciy4jhf5i1w3xOROonaJTDEySiba7Q/KW8+Nb3kpUDjB/oPs2IjmhDmBjJF9buN/gCf2WXB
15rIiGkjNDrbclbGh0fcakTu4/9un0h6JN03Wxdhxajqz6TRYCQO0HUQF4iK0JXLTOsSuVaUg7R4
1jL60iQs7N8T8YSAQRkD8ABoCF1R/RcJCWH6mJUjiKunA2u5p/Xi5fdCdF8axabkfXVDeKOeIMeE
fPjiDU3FzYHmMt3lZZxCZimNb/MT2x3GmS1c+k9N9MXkiGfc8Gzo75Ww02PCZQ6Sw6GBC5HjZD4+
YYkQvERFyCBU5pghk7+z0BkQYrAymbrasWHkVXB4PUF0RCXCH2wKGd4lHOW/Wib1oGyLnZouul4d
64e2wdgB38uIXEo+iLwkjM7DMzg1rCyb2cPANyffc5dufDltkcwh8b8GccC1TMc9rLTOMSzyyJg7
jLGy00wQigsS9ZXPht5Xl4DA11+j9+NYAgGtsQNUvbB2Gg3VgFhcDV95TcJ+pV5vtkvW0OkOzoJ5
d/HOaMG9qzTSvKPtmXR9gCnzN5kkSK1fCj/RHoATdxoIp70G+h+SKSYqpdicXNFI0WII6p6IjK/U
8Svan7/dX2nKN85hW9hkTIlPv+R2FtDDRBG3vLGS5POaAGcBvlNXYyFwg5rGbJGF7okPXCHYSeir
XEdhGBnLFbwlWPm/ZlmSZ5PB9KrnN/uGGhEl2caKUoD05LA7vdAOw+iuD2SQ2T7lhKDyY6FgJyvD
vUH5R62kgr06ysvG+NiyB9ml4hd/0d1tRdKExO3pOjZ1Mz5HdWis3+aNfrP5tT+z8gkBaZU7/PtI
c2V+k0gzeFvfrnglhcsG0y2TvzU9O1uYwJkq0koBdxp/hiVPKSgUjiPwXzhRxXk2DY+f3p5pcNRe
lvK5Z+Pqbtej3zAfF0a1OJ9WIj9IlA8SNdxgc1jzIQg9iKINA7gJM++HCZCX1JP5HBzhUKzc9dDT
5EF1Pa4Y/E0Svpu5XJeAbzfpBcceXWdaU6K2DQT6jbLloGIIalDbFbttLOneVg4T2ccpyE1F4erO
cDHXb38gOVILLOMRcfe8Bg4FIjUBok3qTwPZXAHJlR4ive0++oHPfDHZYkSEWt74fHark/Y4dooU
LYLsJe+YgLlwilzs/3A+FTY9GC5JjlkMtN0PaqvrF+362scSoY/Dkak/hvRBE3S1LwzgmTwhvKcE
GI2c2130Tl2ne07yWg4m9qJPV6hkT2schGm/cClhqCF50xmKCj5ZFHfFwh086fSvmau9qhuuraeL
YJVtcQ2x4gqCbF9GrU+7OAnduaw12/zsab2tnnmrdZ2x13B8kqWVdu7N8zpK6yitVmrLIuZJnyhG
gvKYI8o9JaIpv1qEJZFSCMSOU0K8ckP7XLJoh+VoCD2viLR5EaCj8RQl2KtmGh4+7Jwtfo3xMtl/
JJANiNxuyHa8eR15xwyp9Hwr4JOuax49f/VP4Yt4fkz7lz3ZFAR8ciKatRtD2eoWgm678KhJ6jn6
7A+/neISIunuZHV3+jl/24u2krH6tJp63ed1YriTwitqJu4zRiRGOXpj63zhnlp/UICcQ3joiT1h
uDgmoK1GMRMhO9lLZ428Obp1nNgYjVLj8mP+2s0CWvwBmctraCKLFYv4/zIMO44WRe0pRm8HQ7SB
tzR9n8ju+SnZQjhaSw8Kll89WqeaXPoSEEvssw6AU9hkKlzewGKNkVWNVR2Qude9j7qiX6rmfBaQ
UfyjvAsOWXUv8wlNJ1Of0TmbIjIsckVE4TtbvsHGmYLbtd3wCNlkYEYh9GXXD+9cSrhV7m93KygT
TLpfCh1WpIKIVdasto7J6cniRMe20Xca3TRKnPEPXsPxkjWIfSAVZupzcMyrdF9+0qvZrTAoi7gt
h8FxZAIzEIbFd/qTRnFAB4RyePO6SKhJNOMrcFCo4zJ0BHqDgO+vibdeslTRKYYVt1aLaM/GfSVN
nEXtcMrx1BsGrsWdncE5+HpyxpimJBWE9GnjR9L+Tf9047SUCCPl7x9C4/p/hrAxjEqJwXDLPiuW
zvHPPpW9fnouPzHRhd7Yg4heNlY43gaURUXQkAy/BYX5L7F5J9YnjJoXa5oLwnS14OwWXJEj6iSe
70cijmzGuwIm966OK1AYPHBpH3L/G/G4X6Pc+wgZuVIA/Kar3XZvTT1MyAnHE2ZxbL68sWOD3SRo
HAIznG3EhlEyccaAQ2yt4c6JMkLW26NpT+AbtMtvcimZ2Jb6eCpjmma6NVvmI6w7dJjPyObmZEYS
KrR21O7mRXcUurdMMfmxdsJsSV0DVjQWfeIKgEr0AfbA3gOmuFTGV5zuki8e2v/Sdhm0zUA9Ur0q
59UmBV/f3v1Vujt246J1NesjS2bUcDiSXOXbbtpSqTdW+gG1WlkqdG+yLmFgvLFVbHZdz0WQE1Na
xKVswG2fwJeTms/86h3x5tSVgkuO57rYOWWbMIl8gTlwQWhHGJYjqjfLlk0MDd525j7aoIH/OzRh
l7Dh1uv9cfPfswb+IqHZc+FgSFoWSacV1o1B4onq9VVgptLp2bTnM+Yy7L3KFvrAvDckj3WnsXMb
L+9+v8twskHeJq6KCESKi4hWSoMtB/NSXlp7QRpym412B6x78Rr/tUrIUvXz5T4UxG2ZLYyxR8U1
BO2q2GK0GQKSkd7OvGkZAUMlxGik5LRumRdDCkovp1MYJ/MBjBYNwrmcZRFj9lm53zeSjGu2RVCd
Qf/2UMDzFxCCKhdw/i9JD07BKB9flhXxS+XgJnhO15/O1qbEfZaxopAUfJEphfmyg6mW8LScatX0
lf3+XOnS9ypflUW+eL3VFgM5f0KykbnwTjWj17o5DGn+m8kcqE1i7nKB3R4Rvl7HitrsdcY7c7vA
z6MmGGPYqBCdIbOpe+8ITafjUeDEsvxXDfimh6Qg2jfyJyZD2sxvttDEYSgAl5H1WkAeCkR8bpKz
cW+RGBXhsRXW9/jHGHbS7X3tu78fkNtdzabblc/0v/U3o3cbR19bVUNKwl4EThe3rGRG6SU6SELB
KbOXMUH0wpU82qqoYArjdLdCTfCv2yxB/V7xYMo8glzeHvjLCjcIJ+25TpPbmEvhW0ZH9zwLevQU
WXqSsItKGTXKyYYlmwg+3O+YruKAV8deJ3SMyIqCk3M/vsgh0Z1WKG5sfNjIRT80qBN9lgZVeJ3Y
iujCHTLVIx10DtbYxOx66xFQf3P8GsE/8K9ZgdPoCPUeJU6mI8p44c4x2mfonWfffCoS5Z1EO8Jh
a76Euhw36bXwE1OvMWeqKCJIcJWGn9UpTMdsr9AIwV90HQhYmrA61ExtzxGU3DhB4lMwEUyCoAQW
QWAf/lXucByzvZFnSEmVvuY3XfcByLuv3pNEy8bjJ268wISNYR8yPnbveGla6qKO09LFHdVfxTzc
TwIDY2drK3SHLKl5oCIe6aoRP6k8FugbGPlj+oCXEiI+cL7mlugA2SLtS6lkUehbaNM5TiFrGXba
I6zLTr/F447dWKXSjKJxLbI+rJPu/cnt2bqtdkfHJU/c1Mf8w8tYN+BMCJWpy5U2in6Gtx0FDXBL
zSMLNmVTJ6S+9+5QI8pO7phut2qFC1caJXO2f0kQBjGMPZgYXFZ/CQbvd3MITXd1WCWCyWCuky4P
PUecy7rBpaKHt/jc0CzxCU8dLa4V2g9QR09an95ur4BnPiyh4cuJ0gTSSDS+d+dgdUN1ddgBPCbx
wcd5+lmKNSH2yO/KiN5r0u/2fMdkbRr1+40gXuxnCCj2pe5TfGN42M/O3BI98iqeP8z8LE86Tebq
pQ1+eKJC6tNA5b3Ga0W+lLetTsd5ZqN2BQFNOR9hyQAXhfIBWX+EIFKHZsmAgidFbd68PzMWxnET
I2B/G2kHL7mujegizSrFJXsLwPjWGrBuF7rML+LkW7evGGk73Xf8qTEloTWmLx98wQ5C++ugq/GQ
KeArv6LOPjbi2B0XY/pLx4gTC4F+B284GXnwRUFVmVvMcp/G407P+uk3eE9UdpauxE4jGGDB7ClE
A1KXumHrKkrR21CqTTTFKRp2C6ejt6rOf5dp6zVVivzvWr28c9urxdcLc1YH4ETnp1XY/qsqMbOE
cFw3XyMwmd2VsS2e0d32puk6XzG3TcPiR5kzm4NN4So+RWHtf6A8MaSO03yOvlKtZqoI6xChsG9g
mPQOx0CMpnxQfBft1eqYvXubs3fmOM30GJVKLG1BdGijPFahkGMWbxmA14bfLH+imEp2rT9OdLCW
BKx/JJ4tbX0vG4GkMtsTVWpxWwha/kXe6wjS/hqAzvt7538KByVrk7jzPHAxV+gMCqxtfumtMn6Z
vLJFiFlFOzVAibdn/QdAcRbJiFYXiJjblrAe3ESIDJx4ftdN48zGpiVV4QUaqAfZp8RQitMSaE9h
WrBO3vPt2HA8RsF3EjEgDH8I5tsWncTNS2ReJLgf88XS2fyMj5qzitctcK8miXorIF7kJRniOPCC
pkwjIVfoyKoQHRah+t6jP/xX0nY1UYYjaVdC6NtuWJ2ovB4JhWVACDlgpANwDzSu+hBkzO1o6+Fd
rgk6KUfgnAKJNI7G6+GLc/M+ud/U3XjmG3JonTcmllBg/spluKWyPziN71aoaccDcrLPSvHbLSEs
MAFEKdZy63WgIiEb4wYcPCgxYYmRNkAcGidW9/VouT1laoytJBjUKhbVdhkXsST8qzPo/uL6ujmF
PxLDZAsEbDxjCRL6UKJcxOMJ58Zn9F4WbJNcCYOyUmWwbHFwuEy0qEtIisLdUu31hvqurKjU6QOH
E92xQ9xKVIbU4ubKwnm/fwb6I4drlfvZyOAU3ygCNPF2rEP5ngjcq4iOUaCS3VOfgGkL/xPeDfOm
we393kGaSwv3PGhg7Gh4fy7o1xg5424YCzsCE4MfOz1WwUPWfXOGXaG3PQB/dhnHbmQvfXqtrGZB
S42RzmjErX5T22eH3ilopI8a+xqlrIow20/WOwj4dbkWTs5HWwkzxq9I0CPKj8zv615/C1H53W7K
ztrpvj7iIyWBMx5ZdBZFTcAfN3itD0oloNOuzcTIiRczzDnrPz+xjOcJbblfp5arUu0RbEynQEc/
PfN+G86Di44O7NljvBC4G2Oh1XbI2tAf4kr2ocsZY7PIh8OBXBjrckmbpWVxnNUXabSsudCBMbqs
FD9i9+yn8lLkzul38EUPc8hSEgxc06LLEm/RYwQi0T8qqa4jpVV8yofLybVSaZxMOK2ARbwPjQqP
BjgEZ225GLEDLTLcB4ewOVE3S8ZBqhUhce23Bo9xooPy+OsJZaw3hngpp16AIrM2W6rGaZQ8K7lH
dW6IyRXqBThxPbdCjqDly/XQHopbibxwKB1nw3DKx0veNJjrzL7dEqsuC/KKqZk0kYKUiWIIzoVt
+BN1EVl0o3QHVAbzWFm1JZHMvkcmG2Bq6Sc/BIT31gvkvu9khWlrBG01dx99x6XMHTw3Bnf9Yg/k
gENlCuBckxM3bEWjHR2cEWFw9uYcLDrv0iTmMwrvjCvKghojCM99ofmuKOxsU1zIcazRd2zXlthX
4UarTU+9fDJBpDjQssg1ONLJI8yuZyXxnuXcSDzu6n0WyDRx1qOiNVZPA+rqfCziSLzvoge+WwKK
pWTpgwFKD8K5yAlDYrIYl33yDaXZe81nYap99DJRtqwLwC7sJtyr7eKH2SrYK6j4kMIPuYi3DccT
85REBrjpH7d9IOYTOIhTbn+vZTQ9gRTpIAr2CqVfkMrtsIjtsFvrbnbg3u+q+r1GC1tmaPcI1RLa
dBSZ8LY5zgEsSXqDR2e5VDHFdoKjgGih5e/AyEd9AE5HV+xnA77iD7qBWwCg9mv65dAnB5qRKWoe
gvgo1luHf2ec6XFfXTobH71bcUGDnbNMxkrU3eF9Hv/8ebFjwWAST33s7tCH/VlOm8In1/coADE/
HHp2f8uB8AEw+g6cwXi/Ocgn0hni8+9D5QmQ6ssBUxqMETwrAP0vFOYahPLDy+XpoIl5bUmevyLw
8LIePL09AN7VTF82IOMygqBAUZU0FECbhHvkLDwdc3FFJJ2TEXDr6LplJG24CI3sNkz2cYmqwHow
t/WkP6HnE9gMk/fZbjNYbx1gxBVavn018vX2dU7zkRcoQT+23xcBh4CnQUYavMsHei/OeLZ6Vr6Z
WEJNEJxAoTTnM3nVm/2mqGQPuxq84KOoyvdpqiGuW2Jo9gnHeQsD0JL6vl5rb3IMUJmDG/PUTp2P
r5ClEte0FmsvEXCklvA+gyqr4hQLen0rHPF58r8pF1l3bWRgoI5nwt3024iA6K51KpZjX5YlxV3j
6U3/QlSIe6eJ1DHDeymMoJDd8BvjwJWWbO6+dPmy3v6VVnbvBEQun8QOSkjwjmjbcPBfjWpAr9z5
clzsAuZMneQ7xZrJWIcteP0ENqnJmcIkfupht6qMWI/z03JCyTgNdAUqmFW1pwEygIbe3uIiAiwE
NHllYzN2nP37JTWQDHJVyxD3KVuewDOnYuFHUJQ+ApPDQiqN67GoNXc3qq2orDCx2GrWYJW9TJ5d
EP+vHKFnha4r+nUkMSTmatg+L/fhodXy3613ZR14jV86o1JniIUA8tpHSbpLnFj3ndRu6e47Tudt
xjBOVnmbOexS39cIQ+r2MvucQErF3Sqn5NcvfCZP5e5C81EoQFGpbYVAkvJM+0UINqUb3Sp7brlm
iQZJvZ4axaNBmhgXMK0TNQ0FfuAdNR4HlqX61mPLVEYUvBn3XMbC/Fh6+XSOaQeWw16rdXutSg/4
Jz3uznRbrO2v9bveQAT7NNrQb4U4D9sGcOWGJvsCDDNUSDptb0VT+kn7BrKGSWCP9em7iaspP+0b
3ze/QEfkhhiqtqIcf5thU3ITfSCmK1b/EJ1ESvFxZTWgd4vzak8EpP25PDGWS32TdLZis39ga+qv
oJ8aHPhPJCyoQS4PhP7w16gdGTK1FClkkFeuPwqDVUxVq/EeCJH2nbfzCnMYeCkSHAp+Bv6P8ust
SwL7WyDsKloh6ylkMG264N42B/Ot/CJFt4CV8ysUHhkqsB2iQOJiXmDt971zPxo4+HW5JNYJ+1XR
DxUTLz8e7etiqHYD5/un7hTwhlE++hBnOT7exhdhHiEBjvp4Ti82aVqfk2a/kjTTd2N5nhudsf0n
ynxW6pB05b4aaqL08Bk/j+QXEW/+hfRNnwHqMoJIwbRO+y4k1tO/ks+nOf0VzaVHrtiZDfjVqO6s
qkRy8TcTrMM98/X6t5Q3rSXIXXVVLAK3Dud9kiw632m+W3BrtOuhdagxgJt76dC1CJDD4kQsRbeo
q/yvgGx3cmWoZWYd/y6Bf7GFr3PlflDvHg23bPQrzMsTPi7UX3P1iYR6VtLFw9m1XatLmcJj8XJO
g3JtkyegYKLPKeW3jrdU4vDBzfAC65BYL1YiVOQKjrufaNK4xqjPuNzfSeioNYplNgUBTiBAYcq9
h3DOzpVv0oIf0G0HZbXzztwo9g7SPeUfgOS4jzhcleMMZlU+BAmFWkMONfQ7p0Jvcd1EigmYr0UJ
pV/KSBcsoDevIrL9BsIp7wlB9GcEXeF0/z+nCEI2q+mdld/yzxd2P++Pkw88VZG8zbFmhkLu71Qg
0I4iUHNN7X1ndgPaRQbZIZtl84d9rSEGc8fr2yLa6fC/2wITUy13XqacD/5K1+UgQvMnZ+w0k3Wy
V7M3m7PjWryr3bvumSYL/EMOaOKMXZdCqQJHktULFTDqYfsXOJRXR7aUmPuRqoN2xRhsqaaX/oaM
E2tlZoXvajLtwLbwQtoRI1//bmiu/Vgw0ySvG8ZAh7vNJ0I7U4vAeVfSfexoFm3ynRN7Ez5OXad6
B2TcuEUEhaY67ij8iXI3DKeAw/V8VfMpwENzyc7ReRvEvn2cAG2g6ajxFmQtyCfwdDmT2lD3UHkU
hGU+jS/flh11Oeh5r/Zph8mohuhNg4fb4zL1UlYtScBZ6FKBcex+F7whse7bBBiw36Da6RdX7piV
nBpQgIIj1H/x991Z8Y8bl9Pe0KObIFtOcX3N55CO6sDnYs7LLrkmq3QtaF+6VkhxdsXAx39X1MU4
DmyIbObPkVFKHljW5krHALlwZ1CuWlbwsD5qiSiWgpB37TRfulQEYBA18o/F/6tPM4nmOzjkBILD
5jM1u0vtS004iPXoVr5LMNH8p8uQ9uUpNcVVXeYFiiAoQ4RTe62fcUm9GERnhiLP565KtAgWC63b
UNdY9VR0Mn5zuKCtURXRtY8sso7K/M7VTvnQOjTjA0EkIagj2mT3Oe/LKjiDugqhpOTPyaifbErU
QaUlAZgn4IaUXlGD5fF9tdVZnrV/Dr67e0ByG+wrfvE8XjHPBP6gxMePiBcicqbU+F7FdvOUBYXO
Fjf78MX2fDuJ+3JVvO1rLRJgOU/dO3wEp8QiI/JWZdOMboJ+OLOK8yQ9AskiHCP6GpzwBlkTuHhN
gv5fxwsT5bJfxJ+eP7GJ9LHMYsY/b8fIsxoHvLl7v2SsGb4Bm5VlbLZz4okhqhnFdgTjUqJuZCwn
wltrreNhXWJjt7H5qQ4JqIY+T0Pe+DJNXEiOi5EMpVdhmnFaXxATTPVrPrp2CBpMLFyHxJdTDUvW
jQF8iQeEoDfnj58fdXbi1N3Ya3Z71vFuQWVJpNyVx/sUObg9xv+UmG4+CAGlD9Hz38qxG4LmFg1h
LWFDOvmABHRXEzn9Yu7gD9KMG71wSkArwNnLCP7gVl0esF/71X1luzzsL7vZmf341lklUBqiKxvT
4RDSBI/QtBgpA4wXaqC1K1K4k2oTtzY2NhitFaWIjvmMCW5fVVU5jHo6ngW1Gh6Yhfhu/K2WWHi7
ibFdgxmKNQjgJZSRbgyadLOrIFeYTqk0Y9l/W0Vvx2Y/h5x7k0AD81dd46rrpTEv1LyDMWL2Zkkc
5OaVPMDPiV5fVK1CVft0UlTem5/8elAIcLUf0jOorhSnH2w6up+zQLZ+bdev9D0pFpTyZh7evWyb
p348gokvhuR3Yvj0V355rTKgs+nMrJMSblpb32iB7Fv49bkZnTQ2S1JMW0nhVdlTSOKcyq8QUEyN
meQ4jsOo+RIyoFoW8W07QpZpW6ufPnFYjDHdQppEZwvoPCBVacO/9vXBLQpsOFnCMGcZN7nvOiQK
WUwt9pd4Dio53er3O/JQHigWnlY+RGzmEcCLSy9iS368affVXzs6qWBllSoIkDWYdi+0ihbcFsaN
pvU0ohnEcAXB+zNCUJRlnJMTDsWQx1aUU4ByDmmVo6e4ifFcsSChOeh3I+gG6rS0d03VCzOzPOP5
Q6gUAscyDm6oJJR0G09cNAsI/ZuH7xtwOumKJjdIPTT9rl62+LDJO61ot+/TlNeL/+lgwH/WIT13
QVyNQdiikoHyzfSWUV2+Y/0sl5WNMQkstY68RYQExxgvpq1jEYLsblEfQZlSYmCnYBHcGOjefcTQ
CJLdX/tTxgE4kJX7JtMwuaqHYOU5tvjaE3N5kCXNOCxKAlfPnPb11L+NqJjONZ3mHfN+ur7mwwvv
15elh/rtJNy8JKayTANwmCWZET4Hlspaf0yhekd2tOo6nh+5Cxt4XyCl2iDd37jBTmCByssLQOMH
FR8taUG7T+EOvnnp5yF2vfAhvwIWW5WcXwUI+4dm7l3ap1bfFgjKBOv3vf8S5x+9KKXtwq14Vn/G
BYbb1bSTbXjhkH0qNjQoKR/aeXy3bopLSUQYcet+LdwWE9148T5S7TcRTjSQ7V+5TozYHILRj7zU
weZPecpTUanuL54+VxxO9FIek8kg+VpcwfZFfY/0hyDb0i+I4n3p2CgvtXQw6CKNR6EvEcQHKDsO
Bo1dTu3QPNNZdkEENAtd2zxF341gKrDUyEw2IsYrxRoifG3sV97n/PKeqnUyM2rXSOJoRc1DNTg5
R2+TbHHiM5I7yvnIOFkzJ4EfXxuNLNlHW9AvWkWytRW2DDbILmzEf8x7qbP04HAh+/1yMDv4anxV
mklSiDQTYuC+KNhtSD/QbCynjwH7xR6ej9d4wKD8syM1hSzG8u4O3ZDPsMr/ekaa/K5wcxxJLITX
Rpm+BPfrxF0BPMkwWaYkMtAZMBtX5IfbdK9eUZl7owmlIR1GpKoZRBRQj3l+GtS5pfXtv5lKn5Yz
evcOmYsv4Cdt8XwH373ylTlQTwQ2PbsTZjPF51WBMNRhB/VIeb1bSKl94NAAjoTbe8hN5/ZWbYs8
ufOGpPdto++7IjEWoQQElbqq3z0rhcTbpC6dGgpo32JlFaufyjllsOlPWpIyXUVD0u4y35t/uzns
rzb7cno+Oekd5t4BHzdYq47uLATxx71YRVmvd3spyeJkGIKfcPAEt8Lq+LWhDWPWbxsX1zzZ/7m4
ke3NyLXgicyswImeD1o1/S7LrlBo4IEKOHDOjG2icZE/IpPklnOnlt3s+7bYux4bFymuolCLzkpA
LxB+qG67w8CruOPVxq7qnQBGWppRwwwSv+QmDVDTXEpoLIPWu2fU4G0ZqFZnikkURQx+vFpOG6Y1
TCCNN/h1wxklC3MTJ0/beYbSTTe8bjYqd9LYqf2sIdJlg1lE6YCxzbxBexiRhoD92ziAz6tOrEZJ
drgyPYzmtvV1yJJAQaLRtzm+rDvo4ZP4ucehV032CO/Ya2OID7dosOGkkkDD3okJaIaOStKQK1xZ
eBLnyWzVgrcm8Nk55OO5VZUZyoEsRGZHFGL0dVzTUCgn/3xc7wASfiN+xYqf0+bblAcOy4pNJ9K3
FQApsNE1RP2XpbnK9wP9pS0eMKrohWsUsLphkpb6sdci1gov6Vq+BPqYFEboj/JlRXjDKSIbN3Ks
VQmOS6rndIrfEcWVClyTodPLJ30Tz2L2Qi9s4DCefHQN/9/FHCLz6gpRV1MemE5rSYakvhdHEy85
S6xH3SkhEwQh0hQZwg9+ekHF9bBtiaFrfdepO09cx084tTI+QuKjvue4RIIwMskZY+JGyM/G240C
Ku6nusKSZeE7dsycmZnyj3lqnS1PKuKUY3cPXq0faxq84uRIJnh5KbLkqRO8Ln8iMp/JWD7NCK/V
tDbZ6cd0J1M8+7HUD0WzCfDML7tGLBd8ULl4XmEF2u43qIP2S1IsoRlpjVciXwwHJOsfEYDPqtUv
pPc5ZEZBb9GhQs93OolxbcEPAtosCSrOXW1yAorUlGiCQx9luoZVJdXaFJDAh1omy0xI/K/Kl3QN
nKVbdT7PO0ugIsg8S677WoePkTsxadoUPIfEicEGhghqdp9By4sWwPKpJaWsusYCNfkMA2L1L+dp
Ne+a7/Rnf2gJGAxsxC1Jf4wRdrqeho1zEFqLTzxgJTNDWjI32QbrP/Zkr5uvf4zZm3v1wcQKVLXF
ZT71Hcv4lPsLHTPN9xDsDuxDC7U0sH7GAMDvBi29geEsT+wtFK98bb+3qjNQ2iAoahWMGq7lwUa/
qj7gJjg4f23uK9M3pKv+QU24Vn6gcn9VeMA7gUldcAyvoYI+8UN02GgznEGOifpuO25niWSdjLdI
VV26bsMuk+6YqpFQsM9vM9r5XIj6Ix3WdEZV/zucEeHrwXxsyH5dqih4swUl3I7uqLN34dpl5TEf
X473NLyvuCgDH4BXQTDvlkdYS1m9Q4Ef6w1xGzwKpvGfrfOqiNGViHgOu5wsXbs6tnEtCxDg99EO
iesnMo4hyeUp+R5w3WcWbpBRUzdbAF6E7X3j003flcErE7aS/BdtN+rkbU1MPEJC1q+j3k3mlN35
DhSx9QPbssY8zeiUL1VugsAUxtVTuu8NkJe238i7w/Zk3dOitUcFrA35h3dKwsl/Z0LtWum8hgiQ
t94iOb39DFgdBORJIwVh9EszPuSqsH3xlc2udbA1giGVnmjLfU2zI3PlOhyVAseilODnqlzBx6tQ
nnYq5MVJQLGhCYfEtMOMtBjvQrAhmmmHFaPhrasPjQ6jdswOA6q4nd65Nx2/lw2hO03rug5wc0Ck
463FIPzakjg/ZHFj5lAorMpsx1MCFWqSYWx0gO0BudOmkNURwxJoQLSN/35WrJswFPx45NT5tkIX
009ADdG/l+qGgBCp9yWGZLu6uI7izvDKnYyVrhAsLN1HbjDxM89m6YJTpcjXQLcNzl3Z3WW42Jad
xVcq15usWueVeZA1fDqnWv2YsGljm+qWws7UAMdfA7FdxEzW04mswopkqdJUTPkwBEr5trXbkoJi
cSiA3sevQ2gNYT3kzBy46Ac8X2gPEpOkO17GEFmIodGwV3bPLGJqey2EzEq/+MnMGYAiWSdy3er8
LO7nQK0kvrA17eHQMrjGiGYXler4hd1yx1gNM4MHTb1X5cA02L0swr1P5RW1/w04f99NDhEspK/T
RTUzNxJ5bqg7Oig8Ri6xkZl4LjpSnZxEQlqle/kRHmR1UlJpC8mFDh1ukj8K1VHEaEG+nmVNpThI
K1r8HM1wnV+qoEDX0D2QhBp3E9McFxqa2yoCEM4MGWVHSJi8muZSYNaoYTBhdR6DEfE05UbddvYy
f25jeCDuchspH954M1tXvwCH4dRs3HMtfOQeQU8/cL3KusMAlUBz9v3dJyNp+4hVVHx3899AcMVl
3hdVvT6VP8L0B6jD+IGT8sfekrRpQ1clRqSJrJknECtd+dNoCZBicLCkfHUK/5N8L1+rE5QvfsSv
OaxqDc24FuMTNWWg8c3ZSJxVAuUpQKMIzK9pF0tLSJBE29i7TCYaGwTddhJz9AkbP65wPql0YWmJ
nBbZx3XyvS/3oiKm6l5Du/rChIB6pytHZzOK3zD7RYAY7UjECHl+G7qZ6C/p37oXxYlCLbcLay+J
9JVNHLulzxkdLa3xHIFQJ16Y3O+mwSDtD+zVgkEER8tEWC4qdSrmm7ufEw2K/oPgfrn/X3NdbiPb
/2ijK8lkk+PI/RFtkvWZEIoN+ifnmu0n7fxnKqioSt0fv3vtBpxFBRhcHep4ze/2EWpiEcGWaeLg
sJETTVqECkp7jXFLKmcaQfScOrK6Pmc627F9s6czwcrNk3Y8ALUrqCE4Fu761A4aDO5tb07xioX1
2zKP2pEN4+oxGrHEGKE98ZJQpGzZb47PaaPqJO7u2OLzmNQA9ThJGo5dlKhXnqmrGf4E808L6TKS
RlAW0k/jCykFfYgxzCYzhbvQBphUdSa82EJCdurifVspFKwKwn6JMR083XyxgnLsoZwwKD84F4sG
dZXBo+7uHqek9JDJ33puyU05ywoNQeTZqv8nbkWcgIKovd45jfNwgOIbIVr29ZAj9DeIdLwhWc81
rUa9G0tgRKe0+EHyhVu2ZN5c9DRXehotdlWKMdmnOTN6EER7XXCviY7yOC//3LbQqpAaFs1cTHyw
Q/rUhT/jUFxOrTuw9yS9I3dPXqPBmU4rocc167OgljcP9DWTxAnGfC6tPMOT/OfhHqmHK2Nz4yn7
prNEY7B78rINeqfJ4nmGQi1YUMaH9S/iXCRTDTwzgBAtiYEJPvDLLo1x60Mfm9Z3pLA/ZR/ZkvL+
2e+A9mbaEYVDaVP1ft0ITcj+XfVYX+Fz7r5l4H+JC6kgkw+wcso475x/bcb2Ae0STNEVRWjNx481
Py3bALPp817KkB9JpeqdRVqoZhADNIhJbUeD/qadGIWa6IKgnoGZmLVA3hFLWg8Os1+LkNhuwcpQ
+gRszKEisN9cFjxUX3xSoPqm8smwhxm3Parg9vKkmbic2lIO4nFP7sHmA9AA3Qa1rMwMl27G6TYl
OkmcG90V2tpDHWgSy9jRCmuVT/SuvvrXYEbiE+uEmIQWxboj4+j1Umj+UTTYYPhlQ+Xsjw9me8s1
UUUveTOp7UcFz8memfyHjJg+rCqnimz6/YqF+C6j1QHFDwjTgiU98Um6BluBDt33IblU3qawV/kU
/A9HkwRak5GGZZGVAmOC6AQ6MtOXK215Jk7/pnHRwCSSBQ87kfbaxPZ30QOfTX4PWgKmqAF3hznn
MN5oHHTUkW21ldq8LK8nUnjezjYrO86w51tRw6rGy4YF9rKVIYhnjpgyBE3l6c3gsZXM2PcUhTy8
+KqOlNTCb0Gvj6s/d1obwIB+PYEbN4bi6FwsteajpAeV2irffNAfd7BNLWBUf8TdUB6zC23vJk59
pyYO7fGOmQtBJUkO39a+ox78E5veqEi9TqI8WxUY+f2VYt9jJqvRYH1S8Izrd5gPSLuZJS1bX/97
JH2ShITy1FjZz0neX7A1MxN/vpE7f/l31Y58mz/RDn6BqsjxZ/yXfmoPPirAhDIm6UCzfFuWniI9
yyqvhYz7Bqw/tEVgJadMSq/xTq/FjCiYIUfSxXyxXWc0+Kw0KJT/jgVZJA1HJm/aWoNsNNAzwb4P
8bCwVbq3yWW5zm389o94Dvy2kabyaK57buuVv7m+UCTAivFvIuKTyAXQM8v7R6UqbLKyNdsce54+
eml4TRDoPK8Vya7kBZt44g8xfD0WW4yB9uvEQbNYsoWbsAb8bQ7GtzNk0y8B3+J4xCjNxXMiMing
Vt0qC51l4vmdUbXF4Pmse52Ghb5lB3Y0gvz1mNgbs7gFA7UMEicxkIGtSVk/2fQ8KwuoETcrvZZc
yCyE2c+b5MpaZeIGY5dVixUSbY6CvazbxosMPAUNVb8DFlFu0iu14e4PqiFV1SxcbAD1pgwGyxef
MBvSYOhoa4F28p9VMvnQ8umBrLkBZhY5gWg17FVcKUgews2cw1EzDXeaY8E2XwuJQstnwY2kLKDc
Exg1t6OH38Nychhs0r8VwOzqaS6Lv9ldO9Da8cS4v9+ctHQdlbRq6wD9dCWiTM/HZ5zHHRj0ZDHD
ZHTlC3+HKeIg3YXJBxADeU+W13lAwsRljo2k0K2FY+G2QrPDOHpqtgsaO36ZzqlIPfx34f0ntfgY
tyb/JhrgTOgvuKmuhaBLD3YQArTbOtbhYqOAysLGZYww/fS3jADgWTUGMg/CXgyQsiPQX0ydT5yq
IX9bRigtCAVQSH3xHDU6/aWCw9jE52CxVPgEq0oXE/tZ9NIlpWg9N4p34eNy0ZqwV3UYApZ18nKK
ubeh6jWRi/oPLxAUZWNsemAi3OsyUJ6vgc/vsqNkBULx2H4EvvLTTXRc2nKJatlBu0eLHbXM0yuy
QuzhMfUlNa0lGUDZlPgTSYL2ZS+t1Rk8YQR2FGSfKPksXvFpBjKKwnQBnc7FeDZ1oo4yVj8LXgQI
01IeW38SEX4dZs+Yz2QuuwCQKi9seaGwlwxJqpdqtubhvJ3PsARwzcGeVTsGGDrpqrIgSTZD4ysV
2L5HhpxXQHlU5x17oB4yprREOtYGUy9Kl627OPzWTmcxlHAm8mz2OhJ3bdOGoa8pHvUj1ky+NnUt
KgeW18ubVas8NCnk1HyxCN0tsPaXWrkLnGWXMT91Q3KU24VlSKkqySxFTeVgsYy9JKHqFi8TBuyC
V60t+p0k4Xjtu7wn6+KDJtfF4tY8nBgfTcgj11CoRJYB0DOXBplhcza+h8joBL4pDnhRXZ31iQFi
FoIlDiMh8RxlRrJ+fTXFUeyFbG+HZeS+ymcn/mEcfWl0ls5U+f5Ye4SZoewlR9MGhtpPZC/oKzdc
GYKD2IJyBTiknKzKDBkSOaYdXQLHeW0PVzRjb6UeyD1jyGGbx7C/KQ1OVnnyK8Sfl7FODxfxKaFg
qro4M9g78F5A+aCNMF+djIWPykZwxlBm6QAtocuWTDupyMOTaAghlorC7ceR1Lm8Ts5sB6xj/i/9
OTmxO42fWqsBnBa1UfQoshsEunS51Vf7wTz2YMBXvZGcM3AH9KEspQCRHWnEU36ehNJcCiEtuIqd
YLj5zkyH6zef5J6aWMpNG4P3n0kR6PHkaZAIVuDs1gGgRHuwfz32vXAjCB72Z8k5Fd6pKYyJO/pl
02UK7NiaqwbTWaV86tPSkv7szu20VRst7Z1ztdnXeg5y0ceEar45D7XGzT2q92/Ep5dlTeBhkvYJ
tZsUFCMIL35Kvzz54KfxabRV+ss4thzk5PddcUM8pRG9w+ngtuuRDh6/VaAn5hWXlYnvxuc0uR2R
8A7x8dbie/fwN7dqA9N69SHbtQqbLQ0y4ylPGCVBYBIY0ZPpwc/TP1Xp0wfZXWxEBItmycj5fePD
K4WPYHEGprZQiYUZ52YeUlpZh6UAWscbN5T2J50Iebl+7AZMoXZL32ozI9Uh7awhMM/e+xSptSC5
qX7s6+gAaCCAbNX8sXWufrZOfoPby9kKx/tSlrXrGvr9nhN/eJukMbXhiy9uevIUz9T888ITlaBd
1WrI8crUEYSvgweCHSxSfXPsjaOWp7nPrtqN9U6RadecgAAVq5v54j+sdIwwauS0352EDrWET1Ff
ZCKS9kFY0eqmPCBZA8cYZ/JpY5T5dM96piJW5hSoimfPDCrXOR4GqJrACODQJXx5CTZm17ZEV2V8
mo6wZ7alpou7iVgkix6vmPjm/D0YLNM9G8WBfSzOz42erGB0cyRgltuBpJkb2zrEd06ixl7f4IES
fpGr4B7cfwLGmy1jivW/VLBpSkePUT76YOHR+Ok/5ZW1yOyq/ux74ka2pSF1zoPUPmLjhX7bUvQn
mbTHFWSZWqOSeBM9Mssqz3D5HZl2xOtYf4hbhmNrrIofr2+MHi7hLFwQLOxwvSwjFX4/PurQb1ae
mdwmpdGkCVZrwHdaoTL9PZBdgjlvCOrbDyAw6jUwRhVtL4uexLKQe+TDpMlAnnhX/oUTkKPA+iD7
bc/LLLpIzYMGn7TnDoWpp5iFW7GoeIGxg7BNTMxrTD3YQQircR+OmvYHPPucxYOejg7pmIBap7LN
u1Sd1AAocppGe+K5KT/QHNDKOewOPOAV/jtlVNQnov0GYwEYzlk7jnXajJzVUjWaaNoaYgB+f083
9XPedhYR4bkc/k+Fye+0uibKeQwVHw1pQNRGZajlLrebBOl3l4f23y1QNeaU5TaYcStMIh2RdqOr
kRVeIgNnz2F/pAuRCy6X5mYKFvIdyK3K+Pj/nGxE1WbhHbF/8fCZiABSVPRgokVmlXN4sK37kKdC
23I/7kghllUVApRBrLJDPhdLljtmyBl9mS+kdlzzVG4LqlhgUufXsPP6aS/SJfiDW70vyyegcpCf
2B1OWZcMhEnlfRI1opO2QsdNvbrs1rhCDPv19ep3NMJ7zOOjAq261nQ+61YT6Y5NcwjWGNgWxNfO
rYd+mq2XE/FVHgAPs0clf/AAGslgC1ysZLaLU1m5+Zz5Rb43bkb/cStwQTa0Yf2VsjWdcNWEPOi+
gSDjdKbPOQEuqvMx4QNsnAuEkHxzRCXqe8J6KHYlHHWBlbtGhEksv5jY/iU0NrS2EhYHb54MUu33
5xvOaOmIqwcpME5qapdZgCQx5wL3a0rVjG1A022xP1dt/jpYloQW/oT3R4r7qkW1MOAAvs8m0by+
I6EFaa3C4vdgpA+Ceo/jmTcx8icFtnLcTDdzvPqPs75nMQEZf79/DC3XDrVbYMiX0lAH8pyYK8Dw
G7WX+67n8cXUr8oj+Ev7gVgv3ZJw7DtrRD4RCPA8KyWvPXa16rfZLi+BE3z2iND39NpEBCE8ZfcP
G1GbC7dzHBVmyV2Qb2SnpOgqLVBUA7aR+sR6WzzG3ZP7aO82JA9raTLURHmxEUHvT2G4EpgYEQFK
drbfHmUV5ajk6PFaqB+/967ia+iKJ+Sc5nJ9vjhRMJHADDXl9jOiqlvDvDtM8SMDtOwm/ZlJLzjD
sueoyTmMddNC3dEx9YfVOpT/llciDkQgobe55cWds2BFadti+loSLykYRwtnXpzIIiapCtaOuYot
iq2HGD0BWXSYcd9BAii20LhN5kSm7L/sTtn0HluUFjUInw0gds1Alai/Z+WwswJEeG86TVoeDziz
sAt1Nj+xTFIa7oJMOg5ywzGMuyiCACTm6aFLeqXL42Dv1aBm9fd8DZQgyp4s/1T5YKGpPr8+ddih
wAks9GhaOsrygh5rHFFI186esB4JEdndT2MVBJ75RXKiTPXNsCzc/EiyTwNgQJEPAkup1gB72dAm
hZt6LHdMy5uYDEzl3HDv1BPnFkEwvFKhFKPA7VSTI1Z7KlBld1zaLTTFfZZPJ0c/n2cV86bgXse1
u7bssjJPDUaOu5ucQnoyLnXrcDzvmY3CnbQanyS0ksUHyH6W4wOgETf4JUsp2ihP2xd8qCBnGO4/
qXulF2QvOmgSvbyNBOUpopA5EsRvhH6TMeplt3u2ITce9GvCFJd/J2UClmPlmq3VmYjri2P+8IuN
yPsnlUd9vtGkpRZpsDZd6xEeIj4vDb7USgemXHqRQB6RATljWkzOSW+IVeghpwP/29Dq8pVz9h3q
Cll7ewWHHkh8B5gRmAMb8YDFL8GUAWLKYbUSmjSC2O1giNmxr0sJSBmB2/foBXRIFcRxje0NQVoP
8fAO5PKjaZ+ovrkuu1pZGVsx9QYzwqsia6SPlUstEQSxcC5mEMiI14x4Qm1KSR+8trxrQHN4b7CK
I7dtOw4FlCsxjN3j24cznWmwlB8XjbP5/FyWM1EOzefbqyw8kJbKtQhr3JImIuVYM+KvyRkvM+AF
N5YQJalbSor1YrKTlHRFI22cx+lQ6LN3OWn8mBEVgAuWwb7I82/sCzBhvmH8Prvnmz0tJKyoedVI
OXnR9Ko07eL14IGq1rhkhNzzqf1j8T0Y9jEsQm4iL8m99pPjqFJKNk5LzAFc0AI2oGlmDJj0DbAw
eyvvzkmeqnI82/ZamZN7Q5XFLWDnBY+dZXztDKIgcjOAAM0qF3KmZuui1mqSdUycHI5Hm75duDRn
f/FQrNFM0NsGCNdjHLwt2oIK8kjh3WCNhbU7mkaOjTt+MXNVQYK+R/jzjN/r4riVgL6iDAyCWyQo
vN1XFMWj5dn9Enz+Z71Y91iXE8ytxN0h5toaz4jLLinhx7+uicKwpNsVEwuxuaCwmb9qUh2l8hU+
Qo6u1iUzyz92xjfuj1CcK4N9pwzVj7+TgOPRZZnoob4UMb+9xZ0J4s71tkOO/pFlH5uJJqZkqcYA
Z9K1IXtvetWrrl+Rvvfcdq+4c2DXmFHXBbgw+aU4EVEkJhZkPCEFYTdjoN6NtDNJC6jMpvS1fZBx
nB2oprfSFbW7tbTjLB6BnkcXJ3y+DfjySdx0iQlEW/TP4OEJwH1lWjPi4ksJQ+dtLKYnL3+cC22w
xzUHklnYemSo/x6ts/6I6XMsywg4FC6EAxA+y9lSIJqMY7Dr91MDHOZ7GLVHi3X320H57m9em8cS
6kKml5S0IoDD9ZPECPiCsfRDEXsd3dE4GvdSD0ULlqRpYTWqc6FPkyspDKGOau6piD3BIyZmk5ER
RI+97WwHD7oMB4NomczlOM1bB+ZhDudpUW2M4KwYvfPuInOaqgLu4FXRhYRHngjguqtFU4aK6fLD
2XjzdczTvZpfawuhu1g9x+lqPENd+nUpA2w9qgy3F7v2s94kVmzFAiFPgr0VSB1xMORVR1toU3MG
oYBvUe7KKBJvTpvA3wurrRGaiOFl/F3Gy00L2xNkMcFBbVVGmCs06kgGiU2FgObSmpnyV+rik1bD
3BnjLhPcdveRriPeMlrJ/mYWOwXgsvmmVr9trTLzlREje4jvkyA8Nb1f8pZ1cL2PsMClQWzpVNKg
aEn5DiXZkVxnR1mnjdv+GKslTL9J7TDxSDhO2o1CYzbM3DJkR2XqVyN8inwKhVP/3GMq4Bdk1HNj
HwO1utTj+m7Fbu3YnDZ/7P8Vqw+6rx7Iepi9gAnMWv7HlLKjAOBOjNfYgZFcgonm/p/qW6QHyVc+
34yawVQKzEBGetcB5IlRHY38/BlguEyXYZqQYzJ9PvujKVycBwXRXDda7irVPssMSkXNXYZ0IW7j
BKsQ8wfMUOhZi4drNN5ubJj4O3Vl9mMo7q61cjGbUcA+BmeruW1oiuQGspqfOWA2+3MRKTXoGQXA
qGeLi2F8RaTa2ibUSYZzRXv3153O3Q9Qb9DGGSKcShNXevaYKF2vTgzLLR/Y0+R/B2zTlZWOaT+w
Ofhc92FWeEaAcGhGZwTh58cncqFT8UK69UUUoEDtxdHE5NvVzqGCCAJAWIx7kTCbOcsuABgfDMMW
AABkv8Prt5bq1oBrJV1RiZNfYlxrn/oH5r9b8YD8AFq/0PfQNev0FO1xIIHH3mx/xpdUSGnr4JQn
lRpAK+Kph1jJARIR5tNSUZgF1t4POgUFUxZ9NVi8/dD5pqb1JVSxJJ5o3zVotVahxEXDquLT1sLp
eFNi1A59SQw0Lwq62UKDiXyGpYncF+wyLSUflGGTb4i7FWE5LIqtpSgUqmUUiXmMrCJEKzK6tNSE
6Iu8i/AQlmgy0Ys/EI1cM/iI62dlCCce2KNT+RmGLgWuxGeWB+QglmbInzZUvK7MIm/FWiCs9wv6
xL58ug/wMfHelNXxVG4nWWPDCwr/iqvHFpId2xNWq9X///jM5vazIl3b8QOLTgu/rFs5UNd0PJD/
DhIp8+gNE8k8wIzkGOReOzHlXGqB6nBqrHASvqGu10iRxnVGXMevBZT2zNYtxzKW1EwyfwT5LH+9
VGu6vxCVq2nxeIuUuACE6bGdqPS9cR+4oF1hwQ8b72A31ApU+alid5PKhBjl3tmLcHK5z9DRoD9M
8pwNDAP14p/vyW5GSyOe3lyeO5gjy6cvtPGGkGxs4qvIzsvJdH3Lv9NGLFMeZZ9/oTwYEpyiv/6Q
CNKrlVCwB8s/SxUlLF1ZB7jhJCq5FoftzGc4uvamvbZvi37cPbYWdmNAR6OdBmNnU1xQJSrAPIlR
NPJROy2nBFalqH7zyE5liEYGrQz7xWkMtYC7PnYY8lHvDRMImUOrlBatwN0AEQ+73XBmSc1VwX0q
gYtvyopitwSLZcX1cT7W5lASyqce3rdWc0Ye04IrVZaGdFJgh/ZvVh+hBthoghu+Gjh+P9XIK1dd
m1DyijpzoDYCwgRxgZaMRfQcJp+IS5sF+ktDLoL7RxM4Vb+11zyL1Vbw7yFtozeuo57FVQG3/FNj
s2A5nV0DklnR3MkiDsIEP3dILsrDh2yD0JcGyg36g054IqiCweHtlogqWSD0Sd38+h88UwsAezyf
SipE5u9WEmZU/klfaSWZY2YY2dAE1IAydTm3RqPWHTSLLwTDCvH0JEbmpEM69GcZ10so5qo0xVkr
QGLDJiiptxPxpif+WRlZQrc3rwxuxy2Tk9DBSjkK2hFw3gwqWB0pjQEgBzwYvzWtyyyp4/MQ+IuG
dpFjeBfendRuqTfy4hCRlQ9xCAGgkyyj3U7a+ii/F1V8u58zi7omMyGpCweha2M0wIx2SP/BT5za
fQsXg8KQk/aubVLmRezaBkWZgTtZ77vYXVqbvPhhz98LZxrE8CYBnJ7Rc7zi6EUcPxsFsd56C+hV
FD+uLoQzf5uOUmhXACt00Ky8+yfE2ORwAjetrgJDT8glTVRqDwnkB6lujqpd/P+5KMv+kjmIp7mJ
JsqWmpDOU3CCL877o7S4HWDJB1PfSNJYIMj8MdSFDZmT2bw+Waj+XxgYHRKhTUsmEDQaO5Y9+p1a
il6IkwrlrfNdtnvsxYE2+ztlrA59UWT0r4LSPR8SKnyOgVFUM3IQzVx355BOs+boIDj93fL0tJug
rmR/X1OqwD/TXTp71K5ALVt2S7/FZxJEEc2oGFhjzqBL1NnsRYzkDORJQek+SSvqBR6bx5RRjURQ
jVQcBSw1MmUF2aDn7/mKcL+Y+5urjxsugMayM8JpcR/bMAXBzxujq1A8XryZn8wOOHQTaEBsYGbJ
ortcK36JfOez4Mwa0PASP/WxmrFahI/svEhoiM/iHpg7J19netn49tuau5g6AIUP2pBfwoduJikP
5sw7Dp42G6zAAQl8DHo54qpVVbOjna3eT27ah+7I+jWPb+di81fE7gCHf3acBnN9DI2tBo1Cgi/f
Z9RU4GMEKYNmTNhKjbrGrRPoVDUI6Eq2Sf4MShtPh3twsLATNOOwZsZhPJRlY9+0NVTVdOC9jsZQ
BCHWSdG1rVBqhOtKQ3o+ZImIxuQDSAL2gTvX913FOReIVmsq/+LhVBkhAutWMGnJeHeVSZygSKLn
Z++tMyJxbKrCDAbuHK5dxALErcyts9ix9ALrZz6X1F6gsKgZCkemdmEQe6q4uRTOK1CnsWcMNI3p
ZaG2ehpCkpdnB7698cOIpT70QBV3750WLA1WCwmUzzoFiYF70MHavIo4UfGR0NOLBKdGvP8eyOBQ
byQ65L9Nwg8NE0lQ6rOTsh4cQDMunaZqF6WVboNzQnprQrvd3o1IPSdBoVQryAOOb+BtHJCFKoYi
dGPbAVBAm76xc/ey0RiR6r4G6SpBJy82eBdoLMr9poezLgqbf88JyKxIvkkcdpiQF/3DmX2hsmku
dXUXfBKsVAquGhcwuwwSkqHo6XsjysBy66o3YTZ8JpA6aeAK4iOCPYM+VXDhqXrMdqVTQ8OcnBQo
t/aTmpODDfe6CLyUXrgxwT8U7SQJQhXbQtY81JNQrc3hjpP2EzQj01WYcHXuAvJT60ohwUbPiy/m
3jAhhQGqz67y3J2kgmzXiEzfclqDuKbUyFy+m8dWRxRmNQbrw5RcxliyzzVe/wW4REMt3jN99wAt
eHiVkDfZ99yn1HMkib6b3RtnAeo3GHcGpk7zVE5Qv/ZdDFDYGd3oNFkBVkG9Pq8hC6usD1FUL0lC
fssCdP0RaS36ZAZbuAipSNYh0GoJLcgwFcim8CDvdmVZX9FhkxEfs/UKq28wFusQoDurw2jka3rC
ocxIFJAsWKUEi80WuUqGzv33kzktfdzoVAL8/46sBrkMz60lOdEr1G+UJO5BWS/t8e6vAYqNVAnc
KMU7Az7tRDqE+nqnKCXa62LAlxnbBsqgXcMS4eTJXj9Qj4+SAv4RfUo07Y+4elSUVzw6IoyPEXQt
K04zG2TZjh6vznnTIw9JDMWGQd+39kTaW++fDVJxtmcCE5dtW/sRojv2+/Stv4yGsdWvMgTkZGpQ
m0vrZWBuA4Aw4UEluWIt+oPcA2wKUMCg+Shq46wtqs7DMGjKB3rA8XAjaoMykbwltzL4F/tCqSA5
4+P0a/mdw8XryXRn8vOqyxg25M4RPibZ3+BG3bvgcrGHtsYSSTHrUwVCcF5ukmX5c7pkGDWGuGZ4
YNfKa1d/sfaWZOrCZOI8j7s729lKVBGWaLeqO0JlmzwRY2k0yKhSyfUsVkaNBlISc3968h92CoeT
1Filpq6xjW28JJkwDhQb6JxUx9GC1t4OuqN6jgPDHgE6Mtc7g/A1kg6yybJGI+5EPEutPu0jujvr
LB6k7BqFlKWg1Ii8TT9ytmrDhg7r3adzYQFXJOoSo6qW0jnG+3yS5gmiE1nHF0qFvjKAQ6EBERfG
w8GNzgD/EglWJmCN0zP5MCm+ouR3+Kt4KjrjDcJUlrAV8geb7Z+0p/5Pq7haM1qMMXyR6oTKzHvc
4N5UitgXpPeyM7qZeCRUNJgGdVM1s5arIKiML1NC3c8dWNP5v58F89gpko93Vm7ukuL154BE2Uh7
mvUYqG3wqvdFfpU6CHELgNr9WJwhE81g/piK7xk+Qg0dDDhHfp16iMUSS8GSL6kv88KCVdbymIH5
VXhMhfdUl43d5vrS0gXyfYoQIZSZjYHvMpw6zhHABvFFn53WCW/kIxLVQUP4+MbZSnqe2ymiyh3U
MRKuPKnzZrdAHAHG8pPQ1QFpuuOKJDsOV4crUbYLy1cofORVUcVA9gOUKmlK8iziLMw+uHQrmtaU
b79rT4/dTGv4Tt7oELXdc64AX4nU9D/kYFAAo+BnzGB4vdKloxFEqYBcTEoh3AJJZfzdNudLj1r2
/A//vdPGa7m8CWeMKjjBWh+4S5xGNlHXWmvoUS8mfS4k5RsY1GA3MroiR6X72yyPrw8vFnxpf2x8
S77xJezuKmK/lxxJs/KGonHLXiCi3+pY9s8EdF6KtgEUCDCBuO0hN8fh2PdOajoMNpGOmzTdf3N0
K0e4SoOqloFcAJ52Zg3dXQHXm7sppA2IEG5Db0Le/1DFZYWaNgq9mOvFfeEhkywLa1XnH/enYWqn
I6cMVcD6oZzTldh/17U/u+E0bpZp4biAMOAgbceTgrLznoXbHUOrcDB0SQAKFwbLvvpZeLcauJ0C
BP+nLy3krI5gWdlIHKk8luPg+DaiAaQiIoKjYwNJktXUSAnOTm5z06tjgOHgP8cm+L+II5pCYedn
FeINKrdtyzzAcZ646MEbEpa/jH+csFx7Fd9c6JIgCRGiHTjfmhOYWrE3tRm+9edkSXdSKTXHcEG0
ad+M3HPPEAbAtKR5MN2Fd47T2hnp4e1ngPy3J8BJ0LrHks7nnJyQM0Gn7bW/xzqUsyPhzzhFDq+2
ps2M+a7uCBs8R3I49kaMxrekJFb3ZNE1QkZI1VoUgM5t+D7Xd2N2cFba/fSMJUeVlJrjSplAFplt
NNIjKPMLiCbUZAlnkzFJ4OqMjrfWV3x+PpZBWrXx28erSKkhhs0Gaeyaat9rq2LkHx/v30O2cvoV
qX1qRiNI0hTjL6g34q4YRciD1YXrCv3fYYeL5WREYO1NHNke7S6duLIpKtJFk+CjwoV/w10+zZ42
/qdMNPE9uHSw0X8l6dfaJimwh9iwrO5GRsvUcYYUE9Rd6U9G4hg7ymTDCdLUkZK4plP3/IGoTL4+
PaR9qrRo0VP8Kwep/NgVsb5zM27OUAQE6RBk7zjAH2RvxE9Y8lnpg3DGcmkqzU2VDLw0lSp85iIi
t+Jf+nAptD7e+A2YZQUyQ1Br96imkp7CP48S9lZjESzTVxMfxkpshT4A4+DpcLtPykDvM6jI6YMA
TvQKTHttl/v/iMKzIdtgZlY/4a0w4JTppOk5bW38IEstjGrOaeGkYh/pnfWTrl4wOIj6RPg4pYMW
VwaCj0ehYC3QItbtxPjI7VQgN3uUnspGOeOhqsP7rM7TVqbicOf7PJRYbg3i8keZMK5rfBY6tqA8
JnRI06wQygLUug7QIeURbLK6/bLu7704QoPjSZcUzKLPUb/OJW8ui+S551mY+6SF0o0Hzy4kbDId
JNHbRu71v5OHtWUps5hA3p167DUtMmNLyN6EIB1xhJXEtSNz/SYZCvSICTTgYYOJiEC0CD1GJyu8
o5NAsJauU+lVDwDKH0pCToqdbA6O8c0fN3xSf9C00Sk2XanxLQgpUfkY4ok+DVBcfoX6C/bfBWby
eEChy3GJ5Y4l56CkTmLZSzq/19BaqZAnoydSJBEA3DDac0uR86Vp03c4cpQ5ZEV1CIEsyuKVkI4a
brELMgtEq6Z5mF97R8W66E2wrbYF9GtaCtdwefpwEG877nVAaZQVTVunaPnqhWKrGoZ+yRE5JmTD
+DiTsQZqx9cVUcJwpsiy5UX0A94hn3iwF3CZ4qudOpAnHeF9Wb5jewZ+emJ2hA+DDXl9Pq+ArS0z
ZBTLtFlzxc/pL0rQYuImoDtrT7RME/zWrdvV09ODD3jbFa+PrDOT3E8oLHWlI2eyBjpFdpRdJXwZ
+ebXRJJPM1bqHUQycpHGKENxqZxRYlBfln12wMFx0O++5OS7Ud5aviIjUFmuuniDgse+VYTZ+BXk
UUUG+l6DIBzSWm3QpyHL6Ysfh1BYWqwcY89lj4F2DnQYkfVB3sAiRWTvYmQ5RPfjtBmUEOtQ0mah
ZakBilRVU3uDO89j7rqdfCjlTH1M+0dtydPKbUGT+2bmN+BUTeZfcafk0eTaHcY4VBelN/cLEODw
ZCYzMYpttMsrldmMWBCZnOdEZsM9M+yX0iYOWyuhL049Ch++Pmws66N9zpEg273mWZZUDB/ZFcuS
IUEICqplufTOMdg53cxIzXc8iB1RDuMQX1FK2nZkprPMFK9gT5dfl0KKYHxSAI+jhCYkVApcHaQQ
x3xzj7T8pzhYV3oNBCh5GgEgFs5PRGQknNzgTBmTpj2r5UXfihTeeeFL2b0DButgItDPKm+T3eX1
MjTLALGlfFnrjk2cfdeCMyKmmAo/bHWIWk3CPTMpTwbePOrk6gMT56s+VTvnv0F+kjSljSnQPVnI
jsDhw3f++89BXQN3KQRhA2O1crUd8jZsJxwneaTi/KjOVISjzU6cXV078PTOM6ReK88RowBSa1Jd
JIzrRFqppsE9xl4SAJ0QQBqdZSVwWsZ3UgtH6lAhYgAyb3YI9EAtpEm6wXs+bhUTWy/xBW5t1yxK
oQG/fuFUba4aKRo/i2Suz8nm90YnlHEBW3mkvMJ66vo9d7UCiymgfxMx8vONZONQ2gP2sTa3MMjK
vCHf7jxxScT8BTDXCqm2FapG+4zu/I9ZR1ZU/U/kNFxp3SaoqjPOSU8oBYeOBd4WgwGqndWhiLm3
55ct5djm7++zck9t+9QmDDjTQIyDlzIm82MjmXg6BCiXeyGvm6g+m5DJdEkG52fzQ3MUlLdXWidp
z/GeeSqZvMYf7UuZq/wbnpXxheJB1R4O3KVrKOtpOWwqMMB8ISOggFhx3/zkZD3jcqS1Lwu7sO6Y
9zXGtsEFdCRoeGfRdkTCVCG2/nM6Pn5xjs5RTZuzVogqtQgujUgEeFL5H+vBIhckNOBKoDJ2Vgbf
5U3SqGWEGaAYXFR+Pin8MWn8qnUf1yW/mAy8x+HlIK0ZGz6/k9geMOOur+9W/t+ECE1AV/lk4ZAi
nDmKJ+2ef3RX1Sre9GBzUIGUX/dKFtprCa0f1fevuXgMAfiyzJquywkbL4PQhlRps4I1GoouVHn/
GbxxjulK7GfI51N5fZ+tdFa3kH5MNgpisE+GyMArINwXp7bgqwOQD0q1V+CtFWrBzs8RN7zjrJ4g
mYO6pK2dwGcj7VDb0wyF1mHkgHuuWclnc9Z9p3Ggbc7NS+5vnshMhefd+vPMZhaSzPVC6UsIqm2L
j8tY0x573WiJbB+wuTekIFreY57ZqkMiTFCiGH+cArmk/JmgwKd6hRBuUj7Sr/871Gf272/oxwYo
TbhAuYkrJ9TjQcq0zOHagVa4/lnJmuSH6Fjshz5qGATKvd4NWBpRenT2mNPNnG+JPKxmye6mbbAH
hNhNTFXGbIp5XlwQjvlIgOgBxbLMWdtFakILPHOq0neuH/mm+4z1N8vObPLdhBRDjnNNSSUPehOl
2dEJkDwqGAwRJKYxiP1G2P6gXNNX7+QpcmUqB3MIgIR3APPSb8BJeml4aGO4v8h9LqmQmQ3s2d7O
v8lzC0UiDJupnraZcOOkZRrlAfBfhOtHUNe7TT72+rFU+p9IhGVkg4rj1C1ShFPdi0cXg7r5flxt
01y27q4EqBMr0v8nojZJbtdaqt4lwsXnodEyWqx0kV9qONNkCbR6Q0rkSFWUIO8Ggj9YN2ZQaIvC
OAbQccec4Qi9XvtkdToyeW58zsBukZUPuj9o5oH7h88/xsVN8dxXKUw0Yha3XqH/JJgHpcvZk/ww
E0qsv3++XBWS/k8eBHqJEMuzqGF8fZdVLeNkURhLVcrF8SPFdDb4gsdF6wpBNkafgmnL9q303Quh
igKbKdVvVVt09cOjzfMd9l5Ab4mVEKlKVMM30kXkrQA8PpXlT1cDs8leEP7/BPIBnf4CvChC3cSJ
7VfMEiXSqZ+S1QooKUmkSVsxFnSecq6B4enrPbCZW3JO48mKcaK9x0e1WQVJjj3tvum8fzkBlBzJ
3IBeZrxBYBsXI77eD/wLKuh/Wq6BecE5ZW+Iq9NEQkarkkM0TUIknmvJatdWrA57dgBK1MqlcrVQ
1X1L5q1nqDe8LJlEv2tpPmMcda/slshl4YU/1Uke4z2HXBm8i+XiMKbWjKmywCvHXDIs/GnpSsxD
dKWX/2wk0Koz6XTBKI7BdHrGSzvsDWpr42ByI8PGslVNbNs5N6aHVYca4WOvk6mYVW3KIzvzlYE5
OP/BcQv4vUPVwiV/V7dSdjsCk9coH36SwRhD5zUzVVPdjr865s05kVaDc2e32BxfvPOXCE6NMfr0
WFtROaN+1myqdLFk0PqzCtsJ+OC864hcJniWbfJtPox7zzq2m5d+3mvwGhpiOkSq+vxucN5JLYxf
E0U2gO8KXDaH6G2u5V73HQExfkHPBl3R/DsE2C1lR7d6V9DYImOhLpbtCk3kxppDn0FngDBArx78
hrTN+yZaDJ4p97huxwUObEcvYmirARTNPf2DEKd/ogSpwupSBMHRmlfmOIgX9B+Lw1l7wurfjKa0
/1HNqQgUegb2SBFYDNhqXuqaIoQLndHId+ys1U7ASy0vADbQmGRHzfXk+E7OMrqlqZ6+vlCk6AyU
1FRuM4pdYbykgT0/ZlS+/8nmN/Zh9km4R8djEUOWMSLgpb3DWHrQzYNOJ75AaBfR8TfZ9HYhJG6o
7Mm2xx4KI9fPioGJHPlifE2I2XOHbh2oL4W3aU1SwLl5tyTKWHrox/YfSbL/zCzbD2MWreyG6o3d
Pe78EYVhfBWTYyRw5rT2LwIYkUBUDNMZXI69EYqrQDZEze4aykO1Jp326g61qy3Q57QJAAUm71Kr
SMdwEecpQvEGZ//gKN12APDCOW0XdDsS2rwKtrEhb4treOTgGzBd2NR02MDxFq5w9eBXjnTTJBzV
BJbkqql6lrPB/N7sINFnEFSxGTGSZ965m3dJORLFmUsyXOq6eFxw9pFObicHJQDwdXrDjdAW7Y3G
q9rMFkRvgo4qN/5LEEPEWCAdjMUUOz87OqtU789GkG4mzspneWMXMo5/jOFpz5qPzrlaec9BzgRE
klj18RgEg4zoiOoqU84rZX8aePhnNBs5iPXYzCIagY80jhwPLkj8tbRENwnqgtENNuohHawDOi30
9QlYJypoxqKQKHw8MU2ve/s2lnlhiFjT4eur45uKbKbK1oezukyiFEOmUHkpo8Z+ZiMqgjYMo79k
3AVAN1YUYFyPPT2cZbBe8debvX9Ztks1QO1IVzt/2pGVuv4gUeYsm0zBG1FFKkB/QLQMxLmH3sDa
Poc3UoeeApSUU41gMO410DLR52JuKb0s1oV8Ou8ki6rIykagN/WUGBbMalM8C6CHSaynFmjfFxK8
2a5/WIGClT+/tDPJibZ1E1JFg5fCts4KccWh7d+cpZ7ueIh23o6YxFStM+061RfDlXfOByQRsBaQ
IDbMa28rMTF41RA2A4y0Fj7K31mVsZOsczIra86jSYarbLlcLgxgbBrsjhHY38F8uKqMz8SraFoH
5Pu4/IxJzRhdAAf82JDVl/IiozIpPZLCTthwx4W4bq3XZBlQa9FODwVLlC9xE1msxgK7VPxVXJbi
36xGFKXFk9DyCtxE91vPowpoL/LlbtFBcRVz55MqjyZYvgVhotZ1YG5IUIERsovETMgoz0KiV+y9
+yxvxreaS08/MuSyZp6qS172TCAP9dUgYL0KkxH/3Hr4QduWx/Z2lGG5e7+c20pkLIJNVWIJ1ChH
c0MceXuza/l4i0ak/krDQZu3nVH1UNemJgm5wGofrb2mWcg2MBNhLZ9e0CBZKJaXWSQhXGO5DzC9
hfOOnPEbuFcwtmYbBnmPrEt2B7PUNlUomEaOmaRNEFeeFxInAOJJDDFerI4jRnQUcsOd0pN2qTLZ
Xn/5LU7/hhGJEf1WQla1DcCsy0ak1I9/ERxETJ2OBTosNpP+DRjWMRL581Uw4dH+kPgV+8LkSkR0
TYKGap0w3RwHYznvwVI7fgpv5+kmjAlJ/wp6kLy5Y3Mm9Mb8Tvb6lSKVcrVI4mrwEk5HN2UImljh
1FvQ4Wpfr2NWpmM0lyceVBpnFnjF8Uw40aZ0NNIniMxvh3xy1QA+jdSLU0VQ/AHheWqSILXjIq98
uVFRcbGOZik358KeX231QBCGnVPrCvzgplvlhZrw63i+VlOpW0j4DZfedmtE83HG2yIhd1xiHoQ8
ZbqKF6QqpidCTW04A3m0xvUISzVlpBczOqcjDp0iwfX1sEZRdEXgKmIm1/nokpG5kn8IWsid3527
N8+OT4mXXwHOwd4SAqkDE/WHJ1uTlRpogjfQeiXB7woI1H3ngQEg10PXo3eE6heJhs7x8OhdoJ6M
oFBpaF/fRpeNWP60m2g/071C2bTlw63qfHPUm6bJHLJNlf+5AJvF2Gz8P4Y6Ni67hbKzctaR5JyF
W+Hr4jcCDg6iDv9rQreCMXJTTo75XwoEqfPMniROsyXx47JtS6A5i47l0NxVFVLWDt1ody5JyFPx
TNDWmIrRWfmaDNpWyne5daQExsH89m2aw872/sh1iY64o9Rvqje64x16VlZk3DKHGvpN0kFLqBvF
9k9j7gWwPwrwN+iMRTXY7hsRrrhkf7o9eYFS3h47nw619F6RoAjUzcaFp9eixRkt9gFTQfanf6I+
xVJCRAEAAZWwCLERV3gFq9ONEeMTsO6tkEwfYT1d6d6H8sXTyr2mkhabFwvu+HVfj5nkKXHhRF1e
yR0BBW1CHE6nZGYpuX/nIAYWPIQE96F7tbXYpuDMs9gsP9w7AAMv5cKjKw5Nkdhe+X6CQ8aVgOgg
SWXjXOE13vfi1lgI3TrM2ptVq9VWmH3xGAvi7DN8ZHg8qJdT32gl9/Yn9bLKNapBjGhYVw3oOEe4
ZZpU1zLBFg/e+BVMWtjcCuferaX5ycLoWuy7fFVtBISgUTRk2iWoAanClMriCdrhHbF01/V4kZ3O
CTBkYzHl7TB08yaRJUSR8VJCRlFCuINIUGBoP9fS8kaQePu8Q4CXU2JE88je5B6zMir+bpMXL2QG
QjcWA+O0BYqQmEPftr/206c1hTzziqIdR6+fsC71vMvAqHO046XE4V9Z4zvzyvYZPgK8mh3pMfbE
g5DpzLXY4cAIRDnlqfLNNYZb5qSdl6eLjSLGDm6D2vB36MEbaa5ungZpPOqATzgXrkttKoRJWvRQ
2puPh6caIQxS2MHa7/cr63cBAn04T0wAZFEr/oQuA9T/1KaIT800FmVkuQznGW4yM8H/hllk+1dG
gLdUfFd1QTHM+yZaV44+JQ0TaSw2hU8GzYvnry1JKmSIIWzy/oNzu0uyGikR362nClcf62DQwArH
IgiUE53LNtFBDBVBPx7FjzCsW1qlRFXZQGdUVZ/fvm3RcHQEw59AFG3Tt+9lTJFlJCmIU92N+zfS
0+tsIfvOL0n30QUTQ8P+JF5a+0vaRUUlkxOddlOyT1hJA2zAq1I7c4PNMPrTUyon005xByNH5tw3
FnlBvhY5z1/Yn7TvQhaVY9k38Dgucee/XSt39ziYmT7NovLa56E4gHSeKLHYu9SHE8M2C2lBoNk9
yoKuLPYKzYPOm6jcK/AKM3sAsxE4Seq0JyoGGoS3fX/AFtgkR7JcpAGz42PJhBcRwq6/W3/CUdvA
bPJthFyNHcIFuFhTEjOF/X+EZQTyviOc8bHi9Y6moJ3Jt8h/OvRpxxVBeKV8ZghxTQsPCFt6uLJw
MjTMo9gk1DbgZkkBdflVlqa/SzfrhRSoxj8/Fa0Pn+B7O1EypeGcmPGcnTF/V6OM4FJAdPt7D47h
t0QW0RR5Z/SA09wTxzojn5sFoKSxT1h4JUITUVevfy+JJ1gMOn5kMOOcHPARw4Hm+l72n2kOLX4N
F/soP1sX64/XgpYgTJ14YVARcYIYNOKvGdYm+4F+u5xEvMkiuW1p6zyb+5wUYshKhxHGz5FUv+Gp
TUWEf8m/9v4Vel+bgwW7pgTc6OisbMQGAuCKpKK/vA2CPP+mUwfA5z9wioZlTEynI/SjkXTSh28K
mYNJISX3VLDa55222oNoGPnv9h3ESYbV0aL/YPRLQld1uuqi1oSwMgFp5FMzGlb14wOHX2ZUMjQS
MZU1oyH0ak6IoF96Fl/uhTSXISpJPGbDagmkqhL3rkxzGMe5IvEdEBmxPJ5nxW7Tw1sFOh2Tcowq
sRMmS9l+4vblOvFTWVlZ1F6tcnNIxl0PFpZtCTMLdlrZCc2SxKtyfPpKWFR3rJwSUWPo1bsxUi/N
nlRzO3D/BTZoY2kwFRKX35nDakYjBr5nkg8B7dR5vqPdOpV466QyHIr6xayvFRGCUVnoFbs8Ni6c
P/GDCif0a9QyG01X7nSF5qGSvbaQOVydECejKRJB2VWEEiTdh+e4fvg2UvVKbUi+N4Rd43ZR4wJ/
l+pMETpWQiuEZUbz6kErffMiROKykMpLvG4MzpDPzHLWh9JpgONnhEs1JWaifBdZIEtKmJxusgMp
mJKveFP3kaYi1TJUyPsXzMmBtddlBWN4slAuzAAKO4bPNyrIlF4IVMxha8Ywa1VrF9igHYh9MLuf
d5P7ShB0G20Y3OLijv411walmzIoXz0BQ/h53fTkxllBosMLq7mz2Kj+CVM5K2uM4NfiezfudfUb
aitXkeYevsxhUgZgRnbVTfJtA7YO31VGSQ4bvLD+enifqSGxNkrDVF6hnteaGR4EHimB09jgW2rS
ZF6y12qRla2Q+CXp+1LJEitSiBOYQr2OXe6lsZnUt4Sl6o+Zu22aV8RiyB243AZr4+5G0VIRNW9S
viG8ZyFN39DXiBbvUfFlkxQqYgASD4u21dkf+K2yevDxbYSP+moGKdvWynP7rBNMOAiJKVB1/8oL
kjY8nKXvRvr7vzqmyYN6hrnu9KzJvZWVNMzFJrIut4zbXBHIKLM6Fy2bQuX3o0yEoAtSCiRKKJvn
9ghgKsgsWGBLLLRMgPB41oW14RiKUuJiP5ookQ1cGH+jD3XDTUAqWRfIUy0m9cpQ1fCmKsB8QzDl
CeOY6wH/TTUqp1tCnFbNRDf+wVdnthP5iui7u0SJU49Ve7ryW8gvmmL9lA8ixoepwJU2NfvuODln
gzIJopXM5T1/k2qHss+Rh9QBU9jMkf2IIPxFcnWIDvGTHxzORuMU9daSdGAxvxOQV4yt+azdJtFN
OmY4AsC8UTYe47wNFbFX3/3djYgLVB8a2z+TeQy7+NB+oNNIowqx85OVX0NEOCVE0O5ES/WZ7C+a
ISxGcJG2HFMCI7P/R75AUUmPwH0hnu82K6P26BNFDm7geJxfGMT8eW6iaaZwQziDQ5u0KGBNR5oe
jhLkehZyWGLBhoRYZ1V2wYm1zcupVYtw4krw0FoX6P9uEbJbywnWA/l6Jm9QaYwg/NGhBihtpDkW
qsSAW/7ZmADH2Ezb8P16Dhwv3oudpEOFEp1uMQ7YeqP/7oJy8CZenpevQseiuuCkWgszsW9w0t1C
rBfYmwDhlqgnlpOhtKC7A81MG7kVvH9K4S2q29WyBLuv8j8nGInoVyVOFb0fzmkMWxKugt5z/ESt
KRVUghtWLwLEPq/3VnAOF0pt8ByKF5hNUE/NVmYivLRHbWCdkhEeM66V7f06JHOB/te3ikWvL3hf
gUBoC+zO+8AZoIFSTgjCzAoE+OdoFLo5COCMaF0T6hSQ3ACIzBQme/z81EuMmvTJEBYeRJfHPHtV
fB+ppFN6WFt+yXBrGSDqslRgZEsexhCZIAiAuJU2eCeLt5Uwy5fgNvw0kDEfNNsovnFr2Yo5vUMY
jN6UCncaKUouw7iAaiKpYU9wP3RDHXpAtHk1yYphjwLrYAINdv5T2H54aCIocQqvgztr8qs+kenK
AMQ9s07WrwRsb/ezMnv9EtXcdrTWuuOlM9Yn0Ojlc9FrGHKYyv5h8EjUrmT/RDBmIuAuR5kqQ3fy
WTsoRuh6GGXMZOJWWNIBQekmP8S1JDmR4HpNa3x0MpAuSyi5TYL7BveVJK/Hg6mZLYF28JJqfuoO
iP3bqdelrLG3B1JySeFM+7JPS9abtyhZwjgIr5vrvSkNP1r9CcKLpeo1XHUvSjy/LXQ3PZKDkIfA
nh3XRp/u/hLlWxZqckn6Np6KwG4NeQFolB8mgdnZfwyu04JiihhByiO7i5T4W8ra89waiD1WWv8b
XrVJyG1TCVjDSQ2LZwjNbprJWjCma8qtWQmqzZSGgvnrLbSu7UkyLVcsQ1/uaGT5hwNrj9YBvFVk
tDvOJIjV/AV8WigWD6v6wRpHkL08/2vb3gMszg58BxLdsLSczuiqZzLMxh6wcqZgFHwWd2sMOLc6
0rYRNAErMvhn75Z4zDCith4MmlIkaThriCLiP55IGmAD1GDIywdnYp95ZOe67qGuQWIxz2kHKtBr
2atP32ZhOADOOMoPgkOGbsxphE/vGx5gjF9aJ1x0L0hxKCse5/f7FDB2bBcSKmVxQUdIc4BAAnm3
lJ/Luv2i6IJAJWPpvM1yDeVh6QsB45liEQWuavVscxjfLbr7YH/Tr7tasRqj3xRizycG2xwGgrV6
SOjCQz3EI0jOqq9UwV/LI7bdGI5H6zFxE0fZuyjQV6qvEiaKB7SiL8zGVQs0e8Lu6bJGtdPcsMSV
4FtwiS+U9U3P/vBzW2g+u20HRAM5O+dXG8yvmO/fHPhFrSFv4Iaqay0cR0/1v3UV1nkXA/Anvl5K
be9UB9nPktZLi/ySPk1B5hjJVtNq3lCieNSmVrJRgkbXW56AvijQAzfVrrLWiNu5FbD5/U3eUhYl
PfqcipnSXL2Rjt1yj1vfZRK4+KHtzvx3FjwGrpsBzSCB10laLhUDpS7Am1WIYRw2sY5Sgfe9cPJA
T73+el474SK4rEpJbaadtyGsHBJNheVR5h/rgKnX0JALxE8U/vxNUWnIM5q2K2U0ljCvNChk4Azh
agHGuLHnUlTxLXL4gmKtMuDzjClaK4wRM/5SJUS2P8fqM5jtxrSiqmoQFFVe7Kl8afC9JSa0qZ3/
UcnlBsrnd2NfNVM2gz8MpBnww6aRqcrStJdq87ezsumzdzf4c6X6L/rGGET8xSNkadCVvVa8q7w2
zpifQZ4ZmnRcmBIf0HdDVDNZNXvbvIibNmN3ZsJjIc02TZhBZuh7p+4Y8hQI/qxuNFieHjJTWxGQ
JkX0NrfGHh/nbfVTwiM8HuGG4dkvdBVwV2qHS+EdoE4Yg9NNVN22/5I6hVsl15Tu6u0a+0f3/S0K
LxeE4XdMS5GKTeLGR+D3rkCmdHlXOOiEqTezJEjlVrhuXSwE30eKNzFo6j+wWhDmBmjThLfGTxSg
Q4e+dbgYC+TJYby58EIfSElzrL0klcTzp/excYheAVHTUYmH5JNkAkI/7GXnAPuvm6dO3X++Zrsy
k7yv9FFgOKdZW9jQNZfBiYiVOXMCfbnph2WXTiHSGMyY9m+CJbVZNdxygVRaAJrfd5ARZdIHYXO2
h8p8PZsjGeOPmNIy4engGMQl7dsBg6ZluToT/Zgufjnh/MvkUwmE7EoGG8BJXApJq7tmgGFDCeeY
UYPbo10hrBTsKY/9PekeaDKDsh/Wyi7a2k+C7yBWQSBM3xHIfpg534459HHRIBfowceHlmBtHazL
rrZV21BxayQ+27JQOieynS1WIc+ojMX1yOa7Ant/IwYP9wAtBHNOZ0jwzGSJFRiGTI6ZL5Fncf8X
a+kUgumvNaPHs3U/e/OhMTCcov8HM/Npi42lGDBPmS5ggtd6gzjnqLCwi/GZx+aKSGXELgeu/eLc
QY+ctFi9mZw8ScSBOjHw1nYyXPJM07SsEdlz1iVdi3SMiUDHCfPv17zoO9ezwRvv1ix3TChXQVSt
uzfSkMJMf66ZamfwI6dVPsi6wriS6h9kF2V7A4ng7wZC2+X5JbhFPyxbF17FCxGWLAoYfMsjB8ew
hqoUY6z+K2wUJhevTmefUuwy3NQo3A0JYr5jSFo6hKSZ/MDfdAj+YKN9I6pEqaEQtjjMVG3doTgk
koHpKIOntfE75ju3g48JbUFUJz+YmF0JM42ZGZwt6s5oz8oxqlDZN5Tylui9IkW8SPln9aGXsjnf
uey1U/Z7sQN07tCp0vwV5Hfc3vcP3i97Szojy6DSxQnIQgqPCcjKlkqlN8FiQXRT2Dl1kNE3Njg3
3AjpBIqmYaTgdAuQCaT0DqG+pUV64b6ldTXEMidsZ5qQbIW3sSLfl3iB+8m6R1oKLb0nvqg9J6pZ
tekRQrPvB6pNEkQEOC375EkSqcrw29PwnwvlbpBBl6LbyhJ9GNs3eYO5poW78sed3quB1FbYSR2n
v6e9ynAxHvfhowh0Qy63ZnHNuK23oW6EtWvhKqFuk+Y8cRZugcu2TwKxlDOdUKxhZDdxjMIYNRX2
h+lPFohq2FLLV3Xhd5+RttO5+l3c+TMFxIUEuAHNFxw4URBXjRkhiJWhnAjxOHjtvhsqsqY0CNnG
uxzU+NGYvkAn2JsYKD57aKXq6ctif+kfcVoE75EB5ImbPkEnYaDZgeqTN0q6zCaivs96brwIEVnq
IBEyoG+SR5vARz4fV/cPLS+UI/LZvWXEwnQqu7moiK0/N1ncxfcr4TYS4YKA2YD9uoWyR6HKzC4Q
5GYNPtqYrcUvhLWVwHzkjV/zRjx5ZVQmBtjl2qqVdt/eQED9QNMAPi26hSFUiOVzUZXy4iaKSrBr
0W50lu4DogXeQUDsbjprq4N81r8AUnqyWsKbvsgQvOPlUZP+0moSxjHmtDYsZCRh41UqMsg5FkGu
mVO20leKMOlXWOqgV8ekZOPvwMgW1ChSjglylUvg9qu0fJRT0QiRkybne7gDiVOufaCU0eEf+kly
x9XDfUfdzPP+SgR3pkROLoqeGznFFp6X77Bomc4f+A5+8EuErE0jm+tUAiDf5vf8b3naUtoLeMzH
HlQi8ka7DvOWhuH5cXHOc35vRVMPZ4hf8UfEyt5IgQ0Rer4v7l+E4e28+J8U27JYag9kW1rObFyF
OxEdn1hRPE0V8p4IxOZp56kt/lgAxpHUTSg/uJ0FLQwcbMBw7GIWIVLRhJi0koDIw1m0SN1SV1Jw
cp+SP3hvF588xNp5hCl/Kb/31bafZJuje9PG8nNTjH1oUQlRFdayqZ1EyoBfv5wNNpzxdejXdLF6
fbwnaNjw41b3lvuS/+WM6jXCyVvOdGvLwFgEqGdi9jpxo684+OuQF7Ox4uSStoOpu2LTVqI1ALaS
pq4qws/rvTSOrVWtTQrjbEKedP3OgsfFBdIGISRUZ3oawpOKNzCM6mQLVBIcTwpEQ9hjqtlZmjq+
z6dSunJyHsw2vxAeTIea5KoBsJJiQrPnkwRJ2yTHJiA0+F8npecBJt6o5m+KHxlVxm1SmJHZbahV
Xnl08DkZmWPO1KxGZLjHR/C2CwYAx4JM3dpAgHzewnGqKMDII834tsle0wvfp66galAIcR19Z5XB
9nsc+g9ccK86/Q9dzcCMEtIPBy91D5z4eIMd+M/GnG+x6LiyHpAK1/S05raABxAyyNVOgnmSzrG9
ANr3OpNlfwSWFsMz+iy4SmaQNhtXbOd526ZWpRfSmnqtIHnai+322NOYDhC9MlY6Rt4QCJ1l8DHw
Ef7GTYLaRxMPDwWMGVX2qAuo9RIYYHv1r77gckyodl3OJNIAzbc2jBz7hlIyd2VmOOytnLhAz3De
b7ZO1Bd9al79lMfpq0E8zG5+PbhoKZ0rMz6Xl5FYPmIg7BHjZ3+AtMaYHytjFDb9mdmghnIwvDlI
rkMZx961+dP47qg5WUaAPp7fUoCzrMKBjFTqwdeBDz5uPyDHDEx0U6zi4Tw8yu7aJj3V0bbGGzkC
3W63JM+WI3QUL/7cqa7KbHxLTM2JIUlg89MrU0FQ6X7ChO9jomDcBi+Dm3VO2UBMjhUf58XbeLDX
qOvEvAEqHxxcaEwG/QpyPnVfkyZ/bodsdeMDVbhHaQgozOLxRoZdns1dSM2SjA0CmH+RMJWKxtf4
FO023EgAVYHlDWMJPfeDBl6teinIwq+OkKsrmq2pxqQ1CUI0lLyezGhIWGLiUCKEKuwpicAshQOi
pu4SLn7Jk90ZeuIyGmd82BiNUvVFS4rx7yuW7P+WPkELS06+B49TPpQXyO19UHkFuNrhxVA8ufzS
j82ocgUEGEnAROvct8AQH5MkRwNrtygNfle403dPfp1g0pBSXq4A1LYMyMGXVySpg/bVU95R9V6u
lGsLaZf4+0ihD9w29xOddO9o+O19KpMKBYtDcvnqSZ9qwtojfWG/BHsAvVRIH65OWb3MaoOvLuWu
Ke0NMl4D9OiP/zyR2CLWb91SSXbvnmUUnukm8Es4ZHfuB+XK48DuL6L13pG2s2mrpfmffrDK5Jfp
Ebg6qYpbwBD3rlgVoIEIo70EIb+dwVt7DO/GTdFv5rHlRSwDu3Sm/Pd2BwjBMCKJh/qdBjAsmB9H
qIhcudVX05N141eI9SZA/g1gb1nev+4Cr3Ft8tLDSiHZ9amxcfykm1gEmv1QSeTyB4S70WHk3N12
mXy3lvhBcgosiiY0pPgupIM0JgcrcNbIc/16kEHnxVI11BtqHiWhmwElRSd+taDqz32/zZ38uC/5
RiIBvrj9vtPkv56rJ2C1dXgmSSQWo7drIGt6W8scAKEAxL7cQy/1hWXsDBc9gq8AkVgyMdFMzzTI
U6dXR0fWG4gRnY9VwDKHJAeotc54GfOcekip07bfGNqlfaZOVR2S3ncDjubPGSqZA674f/fD4/FN
jvitWckgEGyT3P6nyQLr7elbGNsXkFy8GHG/rSzk2TeJTx5yOHHccSG4aJ8ejfDHXVcJtWF2bOPr
+8B9WzkwfC/EM7JoGHiGAzzWG3CK5U1x4aO0sGutfsyc211yLfNtqRWw+/phm83AK0iX0H76AYSA
k226MGRh94wpbaKPfKMSmpSHeLllAiTL4QhOcFLQOn+tgvUfFaAazCbXxBxd0wF1AGXxeQ2K5FtY
XlLbbnvh9LtFpFgjGzZge40Coz9I9283tD32ce7eDad0jMlK8D8rtJJHKiNVI2DgsEgkAZcEOskO
9Y8MOYnDeLjTzzQOp4T5YQvOqCinKcV+PqmiKY05NXf1XgvO3Qw4Sy0B3qdgfIemgSHk4sCy+qGs
zlJJ6u+aqVtQ3smXrNUAJdfoLWFasLDnvvKJlmtNVJhPlOuM+1pxv4yKhPVsjKcGOw3LXvpUP7fu
hNMJEX2psr4iA9dxZn2ag90UzMCXKrj2e+RM8yySGwiUv47CKiqWMNiAFbgaAqJqoS4c0iIGNDxD
NQoNpKD6VWqDOkM0RM4JhGIReA1kWyO7DJsq1TJGtE6gRncw+nrc/tvDZs1UAQyhsiQTOh6H/3xB
Hw5peEt3gvZw3HTo7estuWUBD2fgpZOlpfgiy7ydslS4Cjq+/zaldExr1/WVJwdYx5FiDYSfoo/d
sXnQrGJJBINDZHOeVECIpOL9v6qX4y88dEQRhqbbOcXCarBpKdjFkKLrGrhZ70dYD2YZ2y8qhF2M
+Syuc6fwN2d5Ws3ffRTBPPe9hUVA6RN4ioxbJB2HCHmD9KunDPvGTJfMM36d6KpKPjLAVO/jjVcu
yDn+NdkRAg5PoGkEyPu9Z18eibV6OfzeldViVPFAckkbISrvQCREF6oN35dslBiyIj64JIx8nOBT
opvqEIkojr4I1iCkG85XeWfxwtNguksJ5KSavznlYndfO70wYEREYBlPFrTvfBOIQlN1SuK2IOY2
xoYN3p+NJe/k73N5VZhzCgGbWY/wk4RW2CKYlSJHSavaJexJTROxjaLnCQrhERGA64A7gQ29Yg5w
FMCmczCmlYHonWfFKBkQs7crcS0RG5/XrtTMxmtnr0fwI15p0cWTWKSLOTZ6PtxNzuIifb72I1t/
ktq8ThYARHDod2jd0OEPEq4lwXOHovTxbjSzG2mjBTExjx3K4pKzCophXYtwb8vPhN0/ayuKU3pR
R6Zt6VHytpXYhjzfDxzJpkm8f+3oj+TSU82u1/N8v7SmniMaNc1RHf6PQOjHhBoKdbU+6xSLpM3w
mLW0nGlCaWh99Ox5Glkxio0Zyv2hA/7NpCYo0PUxpIiczBv84tGsa1yMgYUGA5syovZWMcowNQ+i
VAEjWvKy+zAaSBiz+Jp79hiVH1xUbcg5P2kpbD4MSvTKtkp8xjgf1m4wPZ9pV4eRlXZXqhaQeg01
NcVstk/65jhEl/mfuv9P0E0HKKn0nje6m95Y1AhBCNImet6elVByVHoGBrsKh+PgEF33RIqM+3Tb
cOFrath/wz9K67+dczvh5kFF0NIx+EvVZamx67aJnww8BYGJvYobsrez2b7VZjaFf1DYifqXENCX
gy5PQEi3Ohv2SzbsJzwTdbMMJablvvhJPmZnJkXqau5uduNbi5Orc8SplsAMcaoBAGl6J6EO7KSH
pmx5Y/BhrDhxng1+ivtneFLz85pkFr6nhvMZ372pF5AVcHMOjeqzL+ckXyukk965hokb6EKLoo9N
wwuMY7j/+wULPYeJcFwZ6JcY9Aygkr2lppR3xmFz+5jzdRYvTNXBIQy/B97p024/uJJx0tK5hb4x
PQPUgHkvXA9uspaADEXwDvSRaJz+GxsAVqYIppGbk7SMViU4kfzlp4Ci+eVKGjZp+qotN987a0ww
DWK7DNUdRwk6Ps5mJYYcVx02utTlXZB/2ergXcunyMhavp9lc5E50ogdCBkmYEeTfbSTxGuf3kQl
722FBRZfI2q13ORsiJC+u5gWTRVA+FC8M7qQi82rZxb+A8JjT7gdV/zQQt066fIW05h2vMltA/dG
9Zrlix+LRrQ30+UUHfJ/tSGwt/XLx5fe9pLl3a3DF4ga804uDEpIQWYPQE1vNVNmlfR1p0flNlVG
yt0aQzCtZEUSCLaR1Q3Lu0osI7jhGjHmeEsc8Vmlh5LKuniRA6b1P+K2HvRq5YAM88brc3Ptykhj
GD+6pdtAAWCHr5+fyN5M9fNfeM91xFpomFL4plRVIgJLiDpBTfwbg1TyPSCzNW1gw9rqwGpHDEHD
gIMi4ndU0d87jpelbreag/RmnezfnmjhiR26FjAiaySCoCJpxPPFuRhLkfQ97tdGz94vt2SRc1nO
h3WIcI4qrZ7MbmFRYptqlmoZAueM0E/ZXGzfAi3Pws9VmsVr9h+7VYkGaFdf1JuW1P7qUGPvgzmg
SVZfxJXDawB/arhjRWdWl9aaA3cHq+5IBzyI1L5h3+gpz9Gr59mTO5Hr2D6S4EGROG8z7WcSNDCb
fryjFYM0DW5nkp0NqewZ3bnBC3aJI9hP6QCWUmoMBBsabwlaQ74vpXnSZE1Y3iwkxQB3SPByzmZ6
oUwiZ3+4rMncdBIdmsqvO3Mh/QkmxTvOYIJuvgOrgqOtaRpX9ZjOueUnv7cKGe9qX4/VI1jO1I6A
u8SHMWQPS26t38zq/230yEzfLa12kpKGe1maAcmkQN6iJozYh40o/zGNJneoaFnAiNy9+HYPtQ2n
RBqkg+R1S/Dx7nFUZPNXILsWig27icB0a0Hwk/DzkyD7MknmjvkeuygisgNcRo0qCy9CzKr4Bs/6
1mpW+VE7Ugdtp/rfpITTS1kwrGDyiHxrwiM3nO7FUAvs6hLFWkJF9UAZgsYAz5VO9+7ljI732eyE
sbOfcgQHyE8JkxhTrEZLjmqd0prLHh/hoe/bgYP3+e9GWawmlqIFmrUEM/T4G1EjeRejsEG1kdum
KKcu/SYpdsnvl6kONAAE0iTLdJSELx7oY5JQj9LOgU4TQEtQCJ95Cin3k/lxReNjVIiTSa4sh1Ka
y+LWi+gablnEY+uD2OsUGpz9rs96LMxSLLg1nt+DfeVZDsy/RJb0g9RPN4A75sMkQy21O7fyjbWw
6IGFyXBEZzuo/LhqCFQrCGBPyOQgSGXsDoR7sw0YyCMlvACxC2HpvL4V8uZC8iLq4sSz2qhahXZ9
vxOb/k6UUlLJNMEiKST3WgLNpylnxrtcMEfNn6X2teg1lnJA3HkB1yE6mBe6yXXOSzN9T1aJS70W
cNLVvfKMsxln1s/3wDD03asVTMHSVFSJVRIi/qa6xWv96DMbY1KxtOeE7fy3sASm9uHn3VE0rcUz
vsEfTywf7J0me0jnNbapNvy8o+0BqAJaQkInyj0aFKyFQw8eEApt8Uq3X1kB4KcQ2mI8H5Jf2aUh
GjxN+8TEK3nVNMkn2C0cYlCp3n+T5mZjXx6sTNcjzzC4C4gpScJyibt9eO02bWuWb4mV0k6EYD6C
xJQMoTqiuzPgtJfUTYW7C/7PvLqFqWZHlE9SpJeB4CWhUaS4UFBFrPICBNOsjSFNUlmHBgEGS9gB
8yztjvVRc7O/vKUOR/YL1lugBxHQqtRCSRisDtCzs+DBTNo8wmJ4dAMfBVgca+5/q7lbCUXQofA6
cnjXzERPu51HMCeSz5k5tVbTueMwOG0/qoQ6fzDIznc7YbZiqbk6JgPoyChZiSFZHpI4Xh5STwLE
BtyM/0Od6xjN11br7S5/SvwSHRiY3w+uNMUOf0WA6ZpKmy/azuklQ7JDbCLMnVPJuwHd+2Tlg+zO
KOEY2jhWfVvLNutgxTsL7ZmVOSjyXYFjtzFNJMXTUVWWZozX1ICI/VN5nFZP+whqa/Zcl7zvDqRA
4MWaOimkBfjp9Q1cQdY7gfie9uAdsAQ979a5aXjXKUKtYYBXeOkx77v6wC9bgNKrkFAltZW0+5a1
MRoZsu8mlx8i4Km0VXUVMFFYCuQI62HMhVTJ/isWA101sOQy7nExqSt0f71sduK67bJARCrmbb+x
XX1eSit0wAkOzD73KnjhxPUWaTg83/zg7V+n5xCfeB4gMk+xb3QB4qF5RACCLVMLYi/M+4luJ9yh
ZGTEzdTqkHt7gifWL1DEQWKaIDxu6Ovykng9qbAN0DsA21J7KuMSxOvB7ZEZBow7QigYuSuld9z0
8q0jYfjhUkZgqvbHnzDwORJKHzQ1MNQUOk2oqh9hQYqqG+LTbLa+4bwL0Ls6ojt7zFKZPV6CJJvy
OL+fh4ilscIODXKAuUqudbMgYAiVuJMwQy802Tuufg3m8XMPDov8ReEi3KnrqEmW29jm/FircV+W
reFgFvdG27754aimFoCqGEZ63AEXSOHt4V6sivAfYuA9FqbQQCqIPRuN5kHA73g7UjTPwCiKwxvm
H8LiC5dEEKVM+vSmgdlT3mtGuTHFXJAK9nKBO0zdP8cj0qJoRhgjAhBpuYiiNH+lDINTlHgf/6Dt
kd60TXx+uI44g5FHCubQ8/p9WzoQ24bhp9K7KdqodvZUYyKHwMQEZxSdMrlxQLVJKwo3n7Zmg9yN
B8iNVROc6R7YA/17krgxZhpwB5VdkXUBfnlX4o5BUww1FoC0rpyXHG8TbHHM4vVsWb1GUWmp0uyb
43gg3zK6j21dxZ4tX6m/IKLSsWTA7Dbr1CXpvZFYxuSMw1Q4HZe07HGBUmCuxG3UgMVuDAXvw8ZQ
lKg8GHsQhKhp5q2g02mztTzGWYXNkBp7oDO1TSm+DCg9+2e5KbzogyFtYJsGvMC+zn60JMsjj42X
l33uwYLFangvoEYmnHRY1s96JYhtRWRLw2LkXuT9gAGiSE3D6N1jKZn0jDsv9bmKrRI6+BTGkadD
6LTn/9q0ghlx7IGXcCetCxCBeL7MfPWtT87WW2MjXCbNgChkwUgBj9E+7x0mWlKyLil0qSxQSvQe
P6nVyy9miECD7wpCzvlPY/Pbf5ZrSUot581MH7m2bo6YTOxvnu2j17AeXx21zNWSOW86wYwo4JGX
ni3pSzcZtyVmK3pVl3II6y1RH8W5bwUZUlrKckcDMoxCeBjvUbTXGOgJekHnVWL3fm/cPN1R00Ci
MMF3ye63/iAamH+XoaYl762OG5YSxtstelCIFfgoMuYIYdPs39zEwRTMZsgQo1uNfysBlukxNzbW
ybrpiWe4mWhKV9iFR3bbBgDss93z/g5ciFD500SIWwW71fshW9hFf+btD8VpF3WXXL85zNLCfrrB
U2FeDcO4QLXCRWpd/pePIRZ+FSOBYTaIb9nBtB8ivW6WC5xvv5ESyxvUdya6QneRzmoHyWZ44TMN
Eq0O0EO1j5sW61jRegT5R7Ix1lyMqBuiShsJvjO39y6URXaoni+tYTFzTFMIFFIZKHORLffx/nWw
foEk7/G98q3lTwnASmwpMsl7rbldLKAct1EWY8C/wmIYJEGLgrxU/xUymZN0mGw1UeVotZW6ak3l
hxQWll8Ih0/ii23fJ3OuUU3iYKfnTklFdeFE+q8iU1rNy11M0RTjRECEabVtdfB7SB76rAoH4o1N
HJz8jeXVTBPjSEqTiij0f/GUUvwIjsAHxK+VnuvhFD6v7hIy42nYL4CWujRsQ2t17HqRaJF7DJ8O
e285aHvRvS8XtivDHSjQ6DV/ooMcrjl0PyafwouwXGOlv4iM/DCbTAyu+Zz3IWJTivIEbKTAwinn
ht1tUbr/TKxISIdoA5Tck6+jUeDJK0kJXCzMAO5DNnCk4S2TLxbcu6/s9tn5pL6instLfhnNL+sl
Ldeuo57ENJmAjPJrguig1q4IN1pOrtWC27jVdqhEItJirJ/nVOvp7rqlIaW0VC6eoep2jt1V7D2S
tqn97HtXteOc60HNcz1knXE6eNMOmDgMi+51qPTpMf5BxWxwRKCSRoZAXH8kyx1iy3oY82OP7E15
8CNnNCnA5RU/vjrPtkgxq3TVjnQdBY759oOWpqEm0oj0ya7wOLfMQ7o0xLpFCgs/FJLA0nW3vLWC
0d0Zu/+WGzYNnY/V1e5xS+DsY81Y/9k4dkMm40faLYl33K/q7vZQRteUS9R0GOVnMLTmEvBL2c6y
KN7LZ6zq6vrN4SJaIMG21+CnXRuCuybLFQ3mnSDEKRwFrLKUxhyBUMuqmu0Y9LXkCFLRYoum/eEW
9oHPttswi2hD4CaWV7/mSVGWlx/dQZwlJAJLC8h3JIo2h5mIKy9QQNQhMivYLZoQtpVU6rKZ8iw+
e8oclKbfRcidSPjmdeZI7T+VdsuNUs2cT34mQEJPes2BYhABaTMlQ346nicU0cAfiQxLtwJVFQhG
WL4YOQrbUMpJt5/bmBuZMttTJUevRdEK+6RZK5FvI+kKrW+OBcY3oxzjMJJrk0xR+vdzNfFBDUQH
aiaXUIyrDIgANBczsFgd7PgcWSmKY/G24FJqtCSrtjhIa0U/vW4ByIKGNiXq9AVbFqzE6Ib0aDMb
gmAwtlHhWCUrFsXJw520quj0+JaDZdJU/0/PCJBiej07yOXFq9oHj7mNUwOQmzRFjJnx07mjMmsR
r0jE99gsHFAM5HvJj9CdANAD15prwAZoOxZQJBHa443uz2rtuDBur/1UbQDjRZ86gEsUH2/snUrD
u3Y3p5WTeVOs6b7SyKuY1JWwkolbEigMZ81Fs5lsIBYKLNphNLwi5BiGEicdGD+WVYUfApjC5Q+c
5m7nM7O1MELzdPmmzmSJDR6BAcJ/GWMSB7QooWFXfJ9wTBANZJdqDQ/T7QgdPD0uPYqtgI69AHQz
qPGzFc+EuMh1PWsYL8n/ilKibh5mBnql0eHUsxrTp3P7H4tRgqtsEpSQn4xpxYAscugoImvD6SjM
8lm+r4SdNAd0rtC8F6YLYAuY41SH9ZP6oBfXTBcn+B7JWENefueN9FKlMpjpfmAfrJA7jMHqxcnm
e36o75dHjTxRDKjWJRHrRu/fVT76ze+STjbBsIfC6POZqeROCe2I1caz5NaeKaIPUBNFtqzC/ZPM
pnnahUJgEeIVSwxn+ZGNMJQnLWnRhX83nP1kTm/+Jyyk+o7bHaQB4gFDmm3hgsQ45bbNng2Kb4ir
Ekdfsc3kajz8AGlhsKmcPyNxZTao2kHs8JQGHf1bK1Xj7IGvwKrCZPWQ0AN1vzR9xzubvzogEiOV
Q4RYh9PczOyE7g3US130pE8bBni352bV24TUbiyflwr0CJhgCQnzyB6th6TFnA8vJVGVrtnvbTQc
5EmWB3TEhpvUkMy9JPkoPZ0s+unPiNbKlEQ4lFojNvjqYYCHvaCFH8DPUd8VkRfUv/rE4FTAggHc
fEBbRIiOJoHJ9Wc0f++AQbaqIpIHdAA0Gc6zdQvMu7AiqQgF8OkoMJAGBJKK6LtJ4Ph9Bpe3Nkmw
ZjNYHjh6CR9qCOZAqAsNB7rNCzF/Ord+4bke1GjrIdqNxGsxY/MYgGu5dYZvoeTN+LfbBuf06nR0
MN//0orL5CjicHATsXzCH+BNvp9npDMJLp97dTzDgD/DvP0Vwwu5Q1uAW70LA2DoeyJemlvTuCJW
DiJR383IigUvu0C0AlHo8664Rd/xYbRcNr7RKgcoZCXNQlPt5YOL+NaYSdExKmxbeQfL2yjweVqI
3Z8qxVdfk4VI6erJOgAUnp4I84BIqhwgILd2FD6UvT1avg/uekZWaAsbpdinXKI02IBqe0qrKnyy
A44dnMq9AWqy61Riht6ybkI0kp6wg0V4kyRz09lxA4iXGOcal8M8I+np/BWi2MwLU/Mw5CmiWyTQ
aQ1c48Oso/QQcFJDLvm2UkweV1ycfGzAeruf7V2s3DTusm94re3g/U322nIlcrWkJ2/SoQp7xfvN
l1I5g9ohdetuguqrvgLuZDQFjpXCdnCZMYUvGeeE1MVOLVVdaEOsr/9sDMIlvE+GBry7V6KE3zWJ
yR2zjPekHWtL4a1foeBAkHZ/S4B7Ex0Gfdr7lzTMIlBmaCMaO51hKczmYr4ojL/Rj1jN/10+ENWC
9kYM8zAt8P4apnKIoeW95LplHHZsJk9K70T1coikwGus9JGBorvjSVCfGWTlideM/Fgz+toHuZoL
ooEm3CUo8CRNHiHpSZzSui2pUUZGyobM7hPUiqvPaAphZLZbSoGAwQV9vR1eoFEbS3guuynvJM2e
Oib89fK9z4/XlYWSlZ4wJaBkj867knYC8YwUudUb6ha9Wot8y/yYZwArq2aWuH8C/ss+199HLU2p
DmG8txk4gr24SWvEVpcSl9bRMIoLWplfZcG1oCMHVObsLTj9tL211MwhkXYZ1Sk+Tnp2HQz3aEmu
4LyckqiFYoacJl4vkLQJKTNwM7h0RREoHF63kCM/vTYqyyCSthPnRekqQmN2f0p28cw5N7r/jLF5
b4CEA/ZfYfx+/vUwTccrjg3zZEEsNGORGweD1IkYBD97YdmDEya5bs+BJvXbvbM12OmxUaqrUT9D
L1kBRycPs65S0LzmnGotCsDJLcwVK22/m36828R+ny8juzoWgnisfjQKgpUl7Dj64ACjG+ZXf3OK
QjD+lQtV5mTHr0qq9AqB9i9Kah1pyNArjgCUNmbjpC1AoS0xjGhh+VZ4/ISvLGacf2AQKeJ695WC
jGn6ctY9IKc666UUOuf8Qa0iXribZEpUQVUcgX+kTYjExLKmz9IBSra2cjYtKIGnr6G/j/etSjLe
EMMjcorS2kj7dYSUUzj2IGIvjIc1rnaoT6+oJdHIXqwYZ4RmYZ3+5bVp7iMlY1S6vdvOqNBJf6+5
17P5+CxLbDlYVYMwtMN8ZDRWeGCJdOT47SQc0rEA5y682cRFofmxyJjd6Vx3ZUrnDCep0OBG9gj+
GXn4bpCwqgZ9EqQT64LCMbaHdSjC9atCtAD8KB/+3V+9/M1dhwWGlhecmSOaIZtbKUYd/35Cj7/9
HF+FCRWciat3dTIfWzQrkE8H8HakBZMu3S6PWVo9yo8nkx8aloyn1jkqCGNxtKCrSdRv77exYQ93
ueSXuy9F9jyDCqUiGQ4LiqGhpUEIWe3BjvEgoyI6T4w/0JGYycncVJ/UZHJAaVjHdkqEvPzROR8Y
NIVJPHRW7EMnfr9jHr/IkGjROybr/WI8Q41jvX9o8AQQ7GTcgN04lMkAxBcJa+wPhwAJEOKqmKL6
BPs5UwAk9DKEFVfm2ZCrLpAMWy5Jhx8sR1gZMJbFrVEKuQQAF+8WGjnE3gz8vcx1ngMbWyVfmlSD
yw/bHfjifgx0E/rAQdofq3wZBJzI/G48JOGy4Ta/yGz8dcfK7Knl2hm7BTAl6NLJy13LWMPHyYx1
crcBM3gImz8nHZbQAtGYAAbQw4+pN97B+rxgUbkh/SKUVWKpmcv9lg4koegBLli3d9YJbf0HUQYz
vm5Hyxotd6xxjS+N+r+lyN0GNhs+bWNDLIcIW6mZuAy+pVVWH0eb4+S95mAbgUiFGm6s9/AluwCj
VyTPH7lsIIGt92J0hckl2gLsuDh1HEWSGPL1C0sWxQexPFbMs6jDmAQglVtqmIxa67A59ZbIdPWZ
DR5gjvPg58UBunly7jt29tpBDV36rtCvvsGMF25oS995UJDVBOOEr4rUN43rvLoIsPioDXHiYIdm
a/9LgedxdT1cBXW0Is8VxskJD5SKXmtfypRClnQpenv1qbv1fVV80fEI+41ej/D6mRnhfgsnQ23Z
2+njOXr46fLGJLJbCVS4zrtL785JiEMwi0IGFOgi3zVUWTrUdmTE3s+XSNiMNf5VutRjK/LNAQJt
yKBaEIe7tx0xgGdVDzj8W8s6arbVyIfCGosVnf/paEu1myakDv7nLByaogj94dSRrhJ4UgACanEH
j2n+AP46bOna+Pe/OcvUM8hm5UA5LNbPdXKTiqouBYEEtt5nxIUzlMUKn9E0s81Y/wYyH6V6LGMj
xnx93aj5C60HKsXxug2c8clduZmeDN+9EHKdF0smRZrjB3mvd/Y3aL0kDhheNrr76GMd3fym1JnN
5vLOGEb4h1zrApKuJ7i3PntWRCYeQlhdpJUR/2uHdCe0O4I9CNMIvpTweGUltlSZSqNMYYynEPD4
1iPn1KPK7w5d93iV/mtvm2hn6TZd02efEXyvYd9tQmjCyYIV/mxFXGHHlax0uK7ane6WRvX2oK/m
Nzo1hZ4XBOJWhS/OD9D34aF4rvY9ROswCETlmpWxnPMx276ySBei4LlWDRC4RNL2Kh+sW7GEeGCz
Uap8La3YVXPzid8ZdJ2WOo11jL5fwi0fs2g+TH/3/mVw9RTyGeLHSq6d7rM6Mj3Gg9z+5oOA66FK
O6HfO8I2qJdx4KnO4yjZGODmFW1+i2OUUv8YGltJPW7oygEaxwGURUC3+MELQACzSfuiCB9mcvdk
Lm6theSL3AFlchEfAp8Jwa6xag8euVd2HeUdiXC468BvkjV5liKyw9E20s2eSP/kQKjngGMummSM
Kn9pGaTyTQV3aPle/6RfA00SpTdi9rPkIkpRpzOGXKsxZVr1T4wDCNwfg3ImzAVXvEMuOeaKbpN1
z+rqijS6n9KY4kkeGMscDGTOFT05k9j3pslqo+GNlXEErCmVSM4RYlVeQfvulSNT8EVRkarQIezk
Q/SMUB2PVJqq8gTOCIxBEZAtog89MgLvZkQd1EFgxOZkC4B6zVcsEComSxOiYoPlvyhVPAGf6SQK
zQQPL1MSoHAf+eao/FB4hd1QuXoC60uwP05rxE1/3G61ASc76P7bGHyZoC/jQT/iFxwdY9KrulRA
TcSCwTWe6Tr0s8WcSbsQzo8pSN7uHJ79r9lHBGEkeQujOZn6mKO8O9LsUHP/t0DR7AMxOP5LXqcG
kzgMdSFNxryMDvlwKF615aIgIzYyBFFmFNKhDxCHJlKJu/GI/jgxNFvzUO5hKQ/5xKko59z/IBRQ
74PdvQtxqKMtV51igiMMKcTazezoZZtSAJZojA71xz8iXJR1YsiYV5XEO29trbSgodcEcCrd5Cwf
e1XvYthUBO/1V4Q4g8U2BnwRc4Ca1+JCfrz8ZrxjbaxZjicPgaSrKWknM9pTCYhaEeVysf5JAMDP
25t+GB709Y90Z5cuOU6GiHv1ao/LS9jO0r0fodKj0X6Xu7cxZ88nuAj2OjfpnJW+V+ampmWV9jV9
eYp6zZqrXg+3s4lIPG4ewqGVuk7PDRt4MK8H5gAymbL7B17j3pgbhiIQ69aGWJTatjwLISMSxM3l
X0ervjvN+qfxZe5xuuv9yhrLMA80Dj7QIR0TBrIKZrTIGZr/BVFTvqh18BMvw7pMVRMLbBkKn6fB
hNRFuOaOenqDVuGNVOZmTjSek7qbEjwJQenAIIQToZGt9/2N8NoRE9xNzZxmDOUJAsQrh4h3AFUj
RPqB7s5RVNgP9mBwHgmUCVoFxfaZZzVY0dKTJmsJacMIWwiU3mEGNgT9tR0U7fGKzsQC2D3n+Qe0
Bk9Li8le9zY9ER0HKuZ0cDeJyrJZQdqXD70e+NtU4TWgd5ZbXCmDIr6f0Hg0T9EAOdJk/xVu6RrW
ia3t+v6ONiOzX1ZrlxV63AjMaPsebJH1Y7p4v5RoQTnoY+z8gXJSXo6oHXZ3MGPWp3hc85Nougo1
whG9vnBD4eXGWexWQ8pfX/lo7/HvILlfCqn0lpcfa7nHSgQWRrbsxtAaq/dQ0vLX1qyjWuE6Tlng
eg/MXOeVZaUGdgBger+duvFdJSyOioBBf3ka/s/OviaclTMdvelHecNgIWZjjbwNyVnrWqB3nJoe
sF3pfeQMua8RlbWI+u4hHsAwyfhJQhccuhmNnR0wgbkMTD8CAA5nvS7QLlzm0BJv186ST3StiIxy
wgDho9d8DsOts7e7u08zxkF71hwVHF/b+epiGbVuMA2uwd2HsOdtKhhfyUHp2jDMspWRSp9Bq+/D
Z7m7YVM4scr59a2OtxstjQ22I9uRGy9iBWgEwCGRNqq02hNbJOU3mPA0iMftoKfD0BDsNpzgmjsi
iEZJWOPMpjIU1nZlalGxBM2o5LG6mTyXgnofnq3KchOk98lQGJ6i23ck3S1IAk18OY0hHdDKP0uV
mMLRMoxsJ+zG7KuawNJy+o6PhrCt8iCD/995mufhW8YlFd9D1AQjnac0u7sdjLQpwFc9ljS2Y1qK
hT4W0kFB+k/LZaDInuGy3K8z/fX16OqomvyiU9XNSub8xU44gTBRxVoAtkQnY275h/o/UAPelUTh
fQxYW/rdPANczhVrcpz7PkFu3uaNuaXipHXKm2P96xEJoYoJT+VDKsu1Bbtb5JoRqgZO+JmAFyUS
f94e77+7uZgae6szIqi+zpEb3v/3ooF0F0RQM3t/dGXjayw1RPbF+8Oj4T8+MebXR8Ob7xP845Hx
gz4qtTUhVI5y7NChCWgPjyoR1kCE9CBxTldYvJ/f4ALaYDy4UbCE3SaF1XeDx4meIDM0wup291v+
i7zTUrtFky8Pe4UdhEeZWqRKygcqK/8NPX+8HqRYIFPDfzik8YmvTJNuzTxM+jZRT4DFRyaCKRTU
Gab/3LlTB6mAfmsNfUOyPPxLXB+oMMrH7wQyLDuXheCp3wUU6g4u2qDt3/hOohXh1VHUv27b5nv3
f+n0qe9zlsfc5v7pzl/vnPToBaCe76KpHsKmXa4kI7EfhK7K5zQn8mCHYpmoXStbw7whLAOOmH+5
uT/yCfIpSnSWqPxZ2whQTBtn7YSVJwcLWrB10pen2SEAtlAXJVyD5ObqyHBKSHQAljGOwDJWMhNv
bPc7T66mP2gsxawb5+fl24L4x9pqFDbsUsoYlskISdK3Fi+h+7OaMeE6vLv+A5vxFARW1tHovefw
94JiCW1LSdgCDw8K+7ME0VoLrzSL17GksKxnKcRE6N8C/FsMZZhd98Lq8MXq5KHCx3T/mx+DMpaI
bO0yRiB7ncR6dki4rZAKpCo4MODxpPkvITqnvlX2PJEg7EIoMxNurWx55pDhoZTaq8bitkS6lQrV
g7uYgEMkKGs/iFll97vslSMwEgOgUhDO6DreFab4fA66M5jbWDBcrAVn99YRWecJikAOZPpw32mV
C++j5uG4p3LWYdoMStIAqSsQU2v+hz7w+kSphke4RbcytOcsSPkrTz32nO6crs7onpV+sm7yK7za
2LrwB8jdqfVe8VQY/2m2/bsvsNMx0gQNZ5nzcZheumr/SybClJ1fUk6Lg6p8jMslmppJp+bquNWp
oSfQDHU9OsComWz/nYMCgbnFiqVm+s+XtlaBd4jRZ77YA0Juh31OWchW4/T9n6OvSu/3vPIqXLnA
4LoKlZN644/J2X3kpAT+KzkEuQdoTtA/VlFBgtMTTg1xeSCUJ3X8nWARuJtjWptKe2900o94Woqo
fLG3aAKgjt2l1MUmbRnk8fmj2Nw43ZfqZlhUjPqAoAkn/ReRVLb3yt7/bCVYL0fMdvAWn0L/7VLL
1sqnhNuHgl0VCb/t/MB3MkBUHxUQSM2MrrGQOTzayDFkRsqf+VqqwFAjLHvOvxK3flv/aAelgb5O
3PlCzggqZLYeE/lvvKOm95jPKQGY77m/Lv4oX86YkHjVMT7Vf9atPsCOR5QydmtfO7Phd2lV9Yq2
wV5+0ly8TjyOjWl/6xhZNLy4F0b9THgcjButFiy4/a4CGuWao6dVxS66ZQ3b7iG+ORNFYWcIIbv8
RzCKDDTvuMJE9LH9tFio4zyNR+uZMLZp0NX6pERCSYwFhZvvVm4mZcHpRtN5mjscjBLUYzGaqwE+
BuarCsNmM/1VxtrhPsq2vq3ysOkyN4M54L3iph/+7MCcESAHo/Sk2JtPmKKiI+NrPnWUFkRpua6F
79X5TmtMcP8ItnWz9kaYFzrEUKhCJWJbdPbJWAd7gE6rWQByhs0/xNtA5ZRAJLVA+iB1w2kpYeXq
h4ZAPp2KChfXCKtfprITjAzHN757zR7ejakorzrqQOUJ+UBZBRzpJbL/EU/danCry6wlURG3V4O4
GeT1EpdQe2akkqISlaPFS68gFaRwGu/hOXrXTo9e8wVFM+Dy85hkfaAfNEoW/RYQ4C4lBcGcwV58
sSft+JrV2udNcIPsbB5PyzTJi7tO3xOuAqzhXvo5txAA+VzJpL0UwTEcq2JvarrCtKbaJPrybrcD
AwFMgKvbwdE1LaNTOxPVMGISab10EAjH34SMqiBhNLpOiwk1x7Z/mgKNVn4aGMow2cVmHnlhfW5D
tjbT9XBMvU3CmC4s18ob5ZKVxU2D5qdBkysaAF4lTnusLpjyYYnBB0V+E+mZimG89+UkYUgqSmRv
sLAKOMFL7Cn4NlX6Ry3E7Lj3AsvbYWZ+S8AwncXZlGSE49sOG/GhsiUgUHDESBKLXK7MUgDARqxw
bD1dkm6lJPk8gu7xyXGgpn8KRpcEtYZ12dNepSc41oMzfUyaHUw8224ZfajLB5JQk9ENTxUR4YTk
epFx9D6QyuZOcEnz0CMOvVS/TAcm2dp43DDpfIIxyarR/eg2l0598/PCIfMlISqwwndCayBJWNW4
08pZhHyHvqflRumx0sjDtbDvhRZ1PJxirgW8MBsMoSBom7WRZD5o7cnz2kySA00SO/mOjDUbELyj
RyDpnRQNsabO0ewvctTcSOlCuI+AwSOLVE9/25jfsubfa3exQc94oG8KqGJZBFaScsiFbDclvq/j
AmgClttsBdqVLKKfYHiYI0ZNBGaKlkZQRyYHNcG5A5o2nvd/N10RBJMOCS4vLDPkZGtjFVfmZCe0
SDsrHNq4tdUClZQoMJc6KVAhbVM9FOB49FotWxjBECyrLv2aIhPiPgxly0i81u0cKbcxI85+xhTW
7B2CjjqZL3X02jTYDrKlHm4cCJTYwgyvE5T5JPTRqJdBMTmj0vRwINQ+C6QaNyOQoamu0iMm8pg2
n829VUd9hVDgAnMA8s6bGEQS3agPnOhbvGhqOojoKPYLv3R0jQo493lcxsI+dJnIVHZlM2xqzpQu
VXZcn081jqg6uyfcJn3zC+8DYQZpm8yv2VgLZ+qEy2z3TwpJRWaKUmVaqC/D0yiH9kaS0BQ+AQLI
RNs6aObZmB06vtBzpbtO4hCvtbkz0Cdf2nVjhO3FjF3xy7zz1EjPlw/+B7nj6g/pmZykkoJUpUZA
fyG6XN6O9yS4d2333aYHDc0/aSOVzscRZSURiZ++yU1XNWQH5hoJlOgmVdyJyGHXk2VGbTwMfeLW
KOibgnNd3V0h4MVvtP09uUZ5eNFZ9KCHiK7BF/LsfvvpslUl/+LeZrlaXJMgO4HDV5vi49G/URh4
sJ1Sh1bjLR7Qe/8PZ1q+G1WTQraq1GAau9AatbObqlzLOQ2VirhZWPbruKD3NehVBOunvFySSJKt
ErQ8eOP5eJUDwbqrmnxxiMOb691SHyux2HdMK4VPXqsFdbfNfNnkEe7dU/JErKBmaFgZX6cl1UmP
KOdHJwz6NbkADzNe4bxOmb7TW4FsPCheQf21LAyv1BmQ+hOmlNe25HoQG20JAiLP3yON5GSDomHW
8A0ApDLQYC1zeFbRkIBuFoqbRWD1Ixe8iowxU34gyV27bYOXKHJioHHAI7kw0AWp9tBm9l2XzbTe
I09qC+PJwTny7YKSo/DDud6ef00yYT4Z1TqLNe9BOaV94DDz4G8gL4vOIpB4ucnXwQAqc4wGC9DB
iyFdyyD6i9Z0qG2LQoT7QEoUgdQuqLcXMbNduM1HI46RdL6+6AtJovBYQiO+I4zUhdXjgOFmJnZR
71bhtVS7GiNUVaCx7smBxt71O1Nb4QS5NW1PGTDiGwQDQRxhicSYARCp4AiONtfUjsQurT+CNLIl
0C+vUGKNoSboJQunjQdh3+F0ydfZ5y4afq3T3fV72gu1Lkrcvmynkq/ODRmPcIHCCp3Sdmz//UJa
/8GMJiRyGFJqc7EL/2T/4GD4lJevgdalDcivMcUR0UVCaXiIYbUlJ84mZccdO+vR+82jZ/kuzcXI
8koc7eOcUQvjtuwgMtSXtnanx3NLTywR4zpdGtG0uewlSPR2IVSHlqDHcQxopL4VH/FI9D0I8HKE
O/0ZC/vyjjudeaoWHQQ3r7l7F70196chxUKTpuHWZu7uBG6XYzrhdj4is8XhhwTK/62fdQMUHz8z
VDxNyBFHpjlHJdJotLGp0iBI9zFBLLt0i4L9S2ZeWQlZqLrIhpTaJCT0YbNPEyc8xs+B/dkU6zOo
TIXlrp/9PHa26cQN/WVeRHNq3/NfD5yE/H+H8EPmrOkg2nmMPUHoHXjnQk2UZLxxIIj4P4/EbtcZ
7vPfQDU194SBW3iozKnBTvKAm4U39E4GSk8AOBzxS1YomD23Zt44s9ed5wkppc4U/OeyD60Vmc4B
iu3KS4dBhp/2rCAy3XXvnsgrD6HOOcxyzd58YnkkmxirEoDPLelnwhdJ6KNxqESPxKD/osEuamg/
AGc87zAj6si7sAX/HND0ZYtZsX51zFwRK5X8CF2OSqcE1lXaBeCC/8UHiKgIYsaxZ5UdUthNF6c6
5osigJnYAe7p4E42Z+nYkfbKXf5Mx4B1VZNdndRcFk5LFkxSj227PEhaNU0QeYh6wFrf+1yMk82u
4dQvO4H9ep6jreoHzNRF//3v7LsdMfXIONt+DDtk/5QSHbVvQYfEUtBJmzIUtg0dFCGTj77JbxAZ
Rb9JBwz9CNLPNe7+S3Ere+yKP2WYT0JLi7bgqr2B0Tz7FpC9pq1uvUTwQmldkAqJ4q3nIkMzU8kM
DPN7GDDTcMrUS2LcXH3v4tr4EssSHfKtWgtzDekysoJrXSVkK80FGl/Iz3/LFO9sG8OeKzWI2jM4
nwG5nD8By5GIZhU0iVe9u23vpSdjf2yZgfxJ3+7TVua5lmEyTj21HcDRZZHXoeR+5RWgcbog49O5
5kztUxVK0taTV5Smm/UNfW9s0v1AZs/Vi/wUxQfxWKJ0a/l/J6dbEa+JY177u/WL8ILWTqLPi2Un
4L//Nd/U8Jvj70g3RvObcG4Damm69NkIQiCfAbkDccl55spF917KAJ0c2oqCsQBAKNpDZqoNLIAV
YQ7/jIQV+irI5a0KwoXlp9JNa8aCzQdT27xVOAi5j64XcmTDDqDUHdQ2TqZYTwexGPeOYoDs61i+
DGvcuKxQXWZ9J5naOMelwqhu46eU0+a1qPX6f+pW5Zea9zxfjBJMGW3Qgp3qYLElkX0+dtuWucKF
u9CDmlvQFVRUSco8alilkNN1OJtDGRERoKPxi8YhtcLSH9LmdvZy5Uht33kkOCk0aPlDw7lCQoq6
aw2bA0EVvzmxYCbZ6+QJiXSTM7/YwVWCHXh326F3CkVBOJY8XaRa6Wdp5BKHpX80X+7JWGEed7jr
HsRqK/pv8MGVk5qk7SXAEIkdAuGOd23O5UrAJhEpvw9UmtSgsbD6NATGc02eNCvYY6vv1QTKFspN
SyP9w5X25K8bzEYP7hsGL0fYakIG32rfdk/Irj1NMqFLmLmfbYJ0Ka5Fq9WF7I34P8RFYpglbj5R
1frqsX8HMhddEoD5emawtBjId2kLNUkNAnxpsoD2d4Rh1P/MTYTrww1Y7OTkBr3texxaHTIyCYYv
1Adpen6vTthMXH816r188gg/OtBk2I7g8kSIdpuvJbo+u8YcL9KSmkGMdlkYsMwVfQ3e9ZFZIAO2
PrpUnaxAuPTsZezVuMt9xpyRV3Atsfv+RXnHyr725tppaPVQDxofw/ExHeQTHubrYvtwOjY7s+Rm
pNZsJ/fkjMLjo1M5G6g7993pkTs3aEOhxobuRaxAWUIm4Iq4NTh4yFJEVzDiJHYVvmUnIVzJLUJd
Ng/0eYwVsJl9ms9xtPgKyb72zpmSnUoonJCstLemOv5iiwyz1cX8kJ8gPDynKTlvfK2TQheHxICj
MRrZbJM9AHmCVc9Q0DWTOq+jY7//yJLUH6qmu9dcRJiWBm61dJgsxpSzU03d5WSzcFOgZPHT6106
ctG+ZzNmHC9XE3Jgv9fGo2t8bwBkLArc5Fhzm4F+aAF55E9umwvMn5zLFbD0hN8aPcesBWCHKJ6Y
lX58cC0BaPa1OkFE1UT+E+xai6+HC5kKS0s4eHfEmgbn7wq3PKEpysM0bAl1UuvOlQMSYZREe1aV
dmkPe1kiWHb+AYDeIM5bZY3A52baznBJ9XDAcCsgSGRknfmLegTI5tCfEwVanDJbjORJb4p/Glfz
GnqOMV2kLzY+bgV0qrsktYYlIbh/ReOUVofO9CvW73lGkmWmn14QOKOCbndaQHE0x3LuiIO+sjlI
9kMnQz+kJFfQB0w9GBDy+u4g6+I00NJ53WgBLToxLi1mEsIl0UlsEseAanfXQpiEj1FlhX5Mn/iB
130bIj7MPw/wo6b8C+TeJlQsVHEaM1+pEj5krvSikW1PzIkhgGZYLbdxR9UuoLvC6+4d8cuPH97E
mb9jpJvHGROSQoxg2LhwMrUTi0BY19VGYaEBq1MN2sCO0cC7w3zAoVdc2sLSEEv5PA3LoCLzltlC
y6HOM16Og/g7NUZKTVWJxAjlVs6d9pCGlY2Tguom8R+LIBvhWyKyYhKtrNlN0b9z9npBg0PtJYN5
fGjiADjyLZfcoqW93EVYrK0xNEZX+zx0sCjR6NHwbYqaS8vPHIKnMnqMJAGf2S3ZlSOQS2YJC6NF
NtjbistWYDX8ejk8W10Di8COz9U8VN6aTFmY1JOJDjaEahlMFIAFSiKZ/F/E7aav6DjFUsIrBRaJ
I6nTNuJqk/XsV/Sqyb+vr7nOpXe2sHyrMnH+P05HV7nJMwVeKk7+UQKVELeKyiN3JHsMz0COIVzW
+dxXIdtVg1VqG44OBvuD07s6Dl7L2CFHf6d/jX5cpy0k1g3GkaMDa8xMD99b8paiz2o9LaUccqqV
exzl+3mzCtPMq5TJOERr/i+IFN++plByCajHiHmiTDze1brsk1zYY/mS262/L9HoJZAQa01d0879
O72nuswWolQPYp+257Q1BxfO2p8bmo3PtqLd7xerQA0nwnBFPs4ye5PjuKIn+Tjia63HTCN3b87a
i2y7Hs74tMLVG4IM7RGFWm4gxOQ/siKtMiY1dhE8gCE2zXIE5Jb872U+X9rIv6QXTrA6J43PDiOW
DINQJXdrrHqTjoBQqCq+0For/LQ/JnyytIggF7/YeWB3oLzVCTwFfzACv7Qs0Kk41Dhwnt9rHzgw
Gs5Im+6H6tkRYZZxPjTGZvNZtqT07NL4Vdz31Wxo/hRjH0abnw4Fj8tRljHwGeX4QbdR26c2cq65
3l1jQgfPi7j37Ms/mfwaqWix/OtHbJ3h/Ojeh2gkaqBHT9AJSguEjRzkSbMxb2kPRD8LEpaJ3okH
PFvplH4084ZM7R7aAVtn6mX8bYYuTMmsxUxUXsgurbzTyi7Vt88VJciTeXpIc7u0jGAYn5VjCYtv
yideazIPUqRQtTN0s6cxOYFdFmeO/VAhHRZ/R73PfQVUfvlsJIXfgX08BUdAJnQJHDYv9zEd3TL1
foO49m+jPFV5kW04JwYo14N94PEFFX0/A1Fx/7adjHhICPTeAJ8SG5AihEI6PAbbMcRhsgtF85LP
gKKC+CmwV42zlXeDI7xXaKAnz9Dkw4Regvkz2zcJ7tv4bXymutJtnQ1vQtCLRFao2gDrYOzDW0WM
zG4gBm7OcITfcVh6PTWFHzlvAZGcagLi6ANSSsZr2wn1IIC0De/y2v6xDCkrr7UCOpyAT5UmPDtL
uBFiqRT6lIOvQ0khpp7GDGsOMqdK+j5dCMrtd/KvNqMPnnpOc2CV3sFLhTHeSoIt/HMB9lrMcwLA
odiVe8y0W7Qu5uyyGAp0xDVFmUmthtvXIU8svIbxv1gwgZenQrF3jGlYbRcThfPr4HW0F5jV8Qcj
y1Sgd4+FznpogJ3Kx7kWwtYSSQBVy7toFjwc2SB3dw7EEE3HG0qKdaXHvu7O0ZhIYDQpFt4g/MTy
FG1taxZbB0Y8IsbhP2Q6dQnZrb8xKZmDZs1JjUknXG79VZWzO+9IL9YyCLvXKFHJWGPjJAi39FDr
//yJRCoagOl5WzF405PQDjvQpkL8lQEjURVPbMkmt/Os4K4nTF9akbhkAhN49+tk1Bot0Zy/MUNH
a9Rhsnq+QJadhIy5BcBT8KprdihBQo5iSPMzEclQ3mfZoK4XsRsL1OpvzXYwbssUXhCUNq8Shdi5
5wk4MQTObsqagqyjYFbdGlbETcrWJTZaTiP8DmIF9tnY6djk4lNuFo6+grAGuulSwgEOeAKuSa13
sTLy66BEOezRwplQZQqYGpun+B538JhW+et6NeW/Bb7xAs7VOyn7U1/vAwKMecu0qO6e6PiDGCLL
GN/gzFQZxnXGsv10ue8JiVNCGFq3kGUl7v8GDTLFD1OH1w/Ylk9hrpaeI9BYRAs+PBZEiM4Jpbj0
KnacCnNPsbXzij59dKskd3tc47SWFLbzAoAmvuV/PDmDn41OI6VGWPEq8F0mHkXRD6o+WONfqoqv
pVMxV9HftNvFHeQsdAyRG4OQyjsn8ZkFBKyQhk/caZGuRvHUDuFeQSuQ+6+U8Ihy+2imu0Tm1Ks5
O0NhGxoVOXrGcq5QQTF2aTV9q9VcS6JV/YyfX2/yqH/XVbuHcKFwFXPBiA7jKVzgSqsL3jQFoy1b
34IuQnqMoSop45JwHZBCIvmD224EWZCnOFaXBkifOyCbnstuCV4Z14NR0Q6xuA9EY3ldq5pFuKeu
MWRALKRxBr8sV5IMtVFsR1Fye06KdFmyIjS2lNKomfztHDY6RtWwjRPgNR0TEeGrnJr4b6tEv+AM
cZ6M+44RL5C1Dx5lBOHPrkLoGJdkMtSB9g9jKMiUx6XOytR97NSUpAkcN4wUn+V87hvjIHQ78tuh
6qq0haDWjHF0VYrcL15qlb3a86N8v3U+xjyM/hh1s4/ZeIKx6PDY1eFgGGWvoR9KfZLINsSOMpBP
5jEGSF3cb0NfkVz0CMhlTukx/cJRIfUwsOIuPzm2902LhoLFtdBoLcYZ+eCiKurNtoBxSlSAQLEg
MDRX/CUz+g0DwJ5XUApYI+Wg3OTXguZRfDExsXlcShE8xH6t6XsRAuDpH3nv0Zt3Lt4dZM4rRFyb
Pyfu9mbYwqnhBYMbNW+BdSn0W0oHjaSdbm1pDHjd2XhUwXJsiaghbiZO7b5TGlxCYvNhGRbvnVzJ
9NyH5i3he+qUXn6BQHeM8MlN2gqBQA3DeSSxbqECSzH8ivNAvkm1tjopW962p/H7QlrIkfet62HX
Sz3jmqxs0p0airGwYwbo5pLNCj6DVnHc3eoXj+YefcWr/PyJT2IP0b95WPSd6y61weupAg1SzXNV
FSy7Ljwj8rkZIXSZxkZXSGqTMbrC1lMcwkyI4omqubzIoDqKUpM2L6Rtxgf8E5GeYVAkwHs4HVfE
ZGID9MJ+d4WarTG90c6E3ufHGxhGUfWNPBw1RfoMCfc7fkawpgeXNu0EM2uMdNvEDzv5b/nS0WJ6
/NLMRqZdm7aaWX2A4yVzN6tbO8Tgy+Oj3K4UggRP3G0ZggCei0sywqqedi1ZWUZqURMSme1oiCKj
8eRLeoXylmpitj5nloRGdoOJhVg2/BHXOB07yPurX1oQD90xhRBk0+xUXdw5h+FlfgtPZcLPCJNG
Mkbf+kSWzaIiKi9ZI4VxZVE1UBikQHl6KD5BfIoXkqf9+Hg5CyiLX5tHcqg0AyamzSoG/C+iw8sz
9UmBGy9dE6udDQD02BXT6L5hS2fkU+Dqn8GXvJDHH0IzTt1HSBbVJ140QWbCYSMdfKIFSTbIc38U
IF39MI1updI/GObjijbE5VIRts9TRMJ3U+L2tDdS2Rk7Tu+MVt/xm0aiAw4FEYJxyWzzmvHvQhsO
8/AaOxgGevu91KRuVdohsid15Qej1OCBjgsmk3lTeIfWrFPFa3ULbuDJ9p36MosCpbhRwD6W07yV
wqXMAwT8qSOWf2XRdL0yNBInlwGrbUTcvKOiCgISRWbH/sSQaZZYPz1erASG2Ywp+cjotLNe/AYT
IiEg1exZyKyDKB7OXeJhwuvlG2k6O4MwxK5eCfAfe9Hrv1IiDYqJPScfEGr/bspDATOW9FlvOGJs
Pgi4HADQX36JL1LySpI4q3wSLN86Q2uyueCaWzhElCfuurg2RFQj3JK59/KoAdJyDGK5VAoE/I+N
YLpUOnwbxySIHAtRPHFjVBBBEFQ8IYRkqW7T907U4q48aEm8ag0s2Qp6iEbv771zYyj+exdFPdFr
uFk+W7DxsSExzs7oQ/UriJKfT1p2P2av7YlqLFWj/ximyCz3H+66YZTyAe2vjqeJQ0ImndI55rMg
X/ZM1yUCoy93CNQ78hbOdDKn95a0Vi7HS3XZHj1C7Xk3882jbM6SSMLlg2mnz+XyNlmZy7b6CQ9F
Ly5NPzv1QgIpOFPGSo6GZB/Gn5kmTUOUsWzbgIeF4mWIg98Xi/H77HVaAUmCEx1wfdlNj5eJFn0/
EuJ0FyV3eytsSxIduiEZdqeW+M5xxYQZcCmfR5KIPoF7FtY934CT6Ynmq1ig3arm7vjnBKn91LdG
vZsygBa9az8PR+L2/FOy0+5au1GqdlDwqmBhYmNOmCyiz7H/DTjt87zxsI6K0zc7RVTz2CCSZ3XI
rTFTCiFz9bXpBGB0RhaQU+iDXynjSmGYXz50g4J0ZjMaNHV6uKZxdYYwXhoVG5rOyui8SLpZGKoy
exPeP2OS5VfpSfz23ZPS23ye/+QUOSeNkeeR96/jynsq0j5YYA2rGeNNSRDEYvf4e0OpGKRLXGyV
il1nslB2BGX2sc+aNAJdDCkhw7ztOoz5owd7Bb9qziDzR4rZCUo6/8a+zQUjycWXcwJAJVMzxrUs
HhqapEAsYV0a/dgRzIXFVEku/sNd884nSqmkSbftSvtHhciW0Y/ZUipaUgnsqSOkMf5VdT7ntI/y
LZf/fLxUe/nsnGNLmFvj5EhxFTEfVCUaBB+lxcxWyzIuz7Ux6sWtUNiUo3fWt6oYlgC3mcqpINC9
HngXsHk/5sPV/XpjIlht35xw9dua11/cLD3W5mU+u973uSQGR1ulDpZhNPcsESJ/727wIIUh/nNh
cStlFfAF0Hr7mmO7g7qBbvjCbI3CWluAsKFDYgu22mE5j5MKmSa2Xv6Q6bjY8YyVsk1kE1oi1WlI
ihzGvaPj+Uhpd2lUV5SHlc9rXaTs32hnImRBSrDKtDhntolCLQvzcGbne0GEy5A5BsbWa0oocgXA
vwFxd03VW9fGfk4Rj5jwcyW95MfrxAtFQtTvbU1q0CiTYhBPZ02B6FVY/thQ84YBZ7qj6C7g/ve9
RvBOtPLla3JhD0FJEoOQLz9Q70eGGJAvRVRRdV+RoJgmK6WTWnVJKDuyYyuGUxWUn4moxt+kwavy
URGra+aTH2EL8UOHtkOrNKdA9IeM+4RxL3f+4aq5Y7+jFUoBr6IACCyIzMtZ5XHSEWYyzNOTVdSM
EPd+niyz8Jra8z+GS8N45D/W4nL9EINicp4ef0Tx88ti1oqLr+aOTXZvLd8zViaXlFg256eetRks
TVVzbV+SrhGMA4HbtWn47orU92gqdtB0JtjToKeBXSYkibzTNdoZi/Cz/BTi5ArjL5LKsmAgpXyc
23NgPoLVImGz7QmuxiE3aRbI2ydczHLSqc5tQovW9Vc7ksKcaxaeV4i77qyZ8mA3Wsb0prlsgVY4
n/i2F3OeY8tctPMdcKTnP+L6c8U+tS9hVe4zIjzhCZPPKos3PwbQ034372uNrnl/wQ1KDKg30STh
X9eY8KvngckWXB+EEpPcSCI7mAddUmXT2ztmSX8YNHOBrVFEub/AGGl0l3x5Wl1wssLAOZgvKMOn
8Eq6qhEoKbdyrUNlu0/wIHXxjLJzF9p57u3N6+BmX3caXHrIK3BmQr3DUNngbWqwcIk7mzzSCuMM
Rx4/x8Nt8eCUjYaauyzWQIeYZhRRKxnztHglV9CCA6MxRBOYxLNsUQbPYtZj2Iaubh81YqSTPBbs
/xQ7UvAsmznWnSpob0nTteQ+q9B88R4rCUZp9pGxoPmdTcyEyMlzPRv43IKMGIMOQRvowbeAmGOl
WzqI+ljPikNathiyGLrJO4CNaS2JqhpijI5+k1ryEXVCmh99+xAC2MukOFLQLUCXC0NTTCCB8lYc
TBmOGrxctZQdvwYO+26Qq/lAIMo+8XZoDnlQD8j8tIWj1ohkoL0DZTwTws6i/05ENoRukDK6rWBb
Xm1AUUMLjmdMfxizuVbVYeiHcjmRoa50JSRL6gNNAvi9wImgq4WmoK6l6ttfa1WY2pCd/urKNJkt
HlFduL6f0T4rDBOO/E9wq/Q8YVy378we6M5q7WCV+CmtWm7akMvp1zDs3j7mV3KAZpB+E7Wm4xfe
iijwX64D/OnulmEtxhHMu+qykcK+JgpOLwfajH5aR74GZsB0s+e335p+ehxG4UcZRhzE90mOMYSn
Gpj1wUoMV1ARmU6yvh0wcXvFK40fGLxms0aq+L3Rc5OAEhRVsrw5tyw65Hm6L6J+7Tc1jcduICMs
HZtr6FKF3aXkxE7ZJF1nt0E11QgyKStID5rvIEj8qsFwtUbHb5cSxxlG9ya+naIwAC6ReCeuy0oP
HwkFE9llbMuTeOPzQAA2RTyCgdxBfP4pTu42nl0QFtnxFYkwuPKouL9LWKfHEgdDOTVQqtrAV7mf
lIuGElS+JQ5Szq5n0qSxhHeCe0/o8yjCnOUlR1fY7JqF+UQrhf0ZE9MRkLafCQOkVMKEYJqAM2Yn
d+gQY2eJo/+tDmobxbTcXlVCeQAbA6KTZI4v4xHXVtvjY60sy/ktSHRMUIqbiAbr/K8gv34n3+1t
6VzPYF1ndIunPWVhbtqDa4USoXOJpwT2gPoYE/2fuBNzRy4CIKGnQ0PCumXYX0636nb+3suV8Zf4
Wq3beCg/SA45o5UGLJ/vnRvv4QB97p28EEKhbvwaA4npaeMl6nj7tX9EjhJVXS2nHUWHY3cUrAuF
q9z+h36C7ziV4q7aD149IgcWS/C2PYozZ7e4HxBFKD8K/UhpUOdSA31fxduNAD4qu60+mEAvMeNF
YkbWdQqUvBMi3i66Po5MTEjo+Ul7gkauiGTMsUwFi60ZFrExV5Pn1tQsbb98EfKMc5ihHfFolkjG
yzXBj6AhV02V1aHniGLd0vmVsxnvnVBg7EQmtD9Kvk/xh3wQKkuro56Zsj0cweUkT/39SRXmo6kX
ZdkD6uhRfLK2lLIa6/Vdr64tE89an6eoz+1iHlHtIqusMQrNkqToP3PeysakDqEgsab1fTci3kvS
yQ/sqcGqS5p0AUb5z5kmhhFCu0JFg3V8fqbqicL0PE6r+9Dew+HUmq38KHRirMsURBNtipqwK8ec
xK/lVroIbbL6i2PW1HFcWSJeG7oWLqOX0N1lob315pY+qMPtNGVxxHQbc/tfjvx6H6CK8vawio95
+Ta6oJszQhU6MrR7ilEu/v0RfI+lWG8CVKNd3iSihD1gX9Z8lYOph1CNWBZe5c7z6KVsiM9og/XG
cl3Z4UwNxqkLptbCNEce2juJ3EGXwdFpfcCJ36S67C+rG3jLv18m1eDpgcM9+wtGWfSmg15ggqSu
6jM6sj4QBdCvhs1ZsdbY7tuv59eBx+Q/Jb0zYJcGnvQ1rk2sTd0lkojLyKQzn58Lstcm/QKBjiRs
3q8+044gTiK+einduxU3/bIC6oxkJCO+KL6rWF0w2Di5resA7+Q+ozlZImtWVdZcVEibNbitEGNv
VWNJOtHdKgGeANIS6014TxJHcP6MfE5dtWZBPiilChVFAGKS6enMNhBgh4OT+8PMpUXRDkFiArVJ
ISj2M678ESkxjSLrh0nwBJmas7gIR3v6mCCBRGPJQb9MfBJ8BfbiBeyEd4rbXAMKcFkXw8zUG6yi
u34BuELEaC3MHpPywmyv9qEV9mFsVTPhx6sBQRwuYDBMZeqKoqFUXYUVdhdJ861RxYUFZ8SAN59Z
yIFdLnrOnDmltiYDlex1BgJ9G05oDCUEix8chVvVfiVnWaFXqvDP4ORXQ8sU+c/NoXGxIBPCmRbY
CtFMeLEuG5VTdfkKxCH2VFO0344fgM7XREIiPr57P/jtFB6Mh0DQQPZIj4MQTFvc9GbRokBR7dpI
h3Pice6YcHNkikLuWx4gupF8xww5vaB3cl2vFrMoM+7lCe3nhtBez/yPDiQoruAgHh6m/GIKjrwv
Rf/OWOtGF7ha7qkCiNGdlcF2ljA+rJGo4EvXtkBRLd8aCkEAv1Xiijv3cdFkafCBg1UQAngOUshQ
wbmEaUw9q8W2y07zFMcHcYiMgi9k5gOgEO+rk5qTUr9ll4qG3t6NFPQfpKsfYvT/jkguako+ZWGS
LyOWMisc8t3QnyeFoqnz7ZfwPEYu8aXhL/2pYF1UUSSPUid27w1hgj2w8yhrTYERPFVPc1nreqrp
WlWTcELRzDna1V4LnEdzm8JiKh2n3mag1NYROhczdRzRahhC2WN4yZQcDjSxMbnIrG8/bXSQA09Z
2MViGtAJKsy92xkV3Lkmg+lbAxtfbw1OJIDMACcrMJRWkHhRYkBGRFvN/FPqZ7uEEPM0gGeTIg2K
/hQizsxUAEN+lVkEsxcn4YbWxiF5gMIFIskUDEKdEnFqtaJ1gz4AEZb28jNV4nvsqabGM7Jh7d81
OuK5+7WXmcd/oXgM3IbBCGzT3uVSfni1Z8jT6Vsl/WbEcWfNbKqN6sgq5CRoZUj5+lJPs7HWL8z3
e+0nwRYumWtmwYS5tvb/1Xzg8fbaCfG/3zBx6SYO01603SMhnSFrnrwG7cm6eNBuUoaVQF6UwrLM
s2pGSFKG2DMPuN0yqPGh3huIzzqQKg89L9c9nV8otmE0FewTx3XLsxGycfneeav39JCux0wvIDHG
b6zVO8iNzzRQz5PW4Wpc13dzxQdEFOn+4VWIdvM4qoJk1SwV3Qnqpa7MAaJ4/+FVkqjhb4O4spJV
tcUtXcsWTB1W8fIPjQWuR11N0t/zpoDevfZVpFZ1VEuKZE1RfPzX0b4VEP2E4BX3OVeIM0//Q2Cv
eFrkjpCNctzDfxW47/dJ3o7lLKNf+Ej3KwF4bkjnNGDy6m/1vH12oEKDh/Kn0jF48KW0SK+oeyHf
/Owu8OzUE/eYfhT6VdrJCDmUYxbVUSq+0uVecF6NNAMf2JozBWSHGLoV4jpIV3oMTeUZ0WoPjSoW
l68k2EJlSsGeuS7OVETZLWMO9d6foD1yQkjqMEtJ8b5+O2EKRrXZvJAtQROFVfmDvpM3ZvwpC/ZX
1IWmJim8g3TJp4Zuki9Zf+9teBllvENKeMi+L0MfHjt+jCdLH9lC/wkELyDotOaklyIu9FgNMO7I
ifLwIgSkbcKVl1jmAOu3ctf5jFiEzgCyKmFCv8pY5IrOPb/f9zfscUOIY8PVUD7R0GUvIuBO0Ke6
rwxB32zE3FpZOvhO0e797gq27h6cQQE5GC3Wd2tDAxVB42dn7Mq1Ks89+VkASsIsj9QidxwlKbN+
LOohNIyt89HWLSjq7JrzpzRkOqeEikV3AJkvFX9IGnf6Qg0lrXCkxfck9/fDWUs0xDMDKAZ07LCA
7eyKhT3L53SIBgM3JxBDSz9bXd4kz2gDqGImYXXBHc8QOTT7qomNdMunSNqPmJJ+JX3t2RoWj1cV
LoJBO3hGfZVW5j4xchgcb+rbqI6cKnc+iPcu4TM6Zkdmzl+k6nvkqmq/1qWzN1/pL71mMa0ZwWgq
ArlzIiJPk3bLyK0NrpifUwGZKzSsXJL4OULG0yngVzWBMQaFHIwJa2wDG5l9S+8hQm0EnibUEeHu
vM9pF+EPNGyGQYV8Tw9ep4wOGmZ2zEtZXDJ86zqcy4mag0EDTk2Di929ajgMsBVZl72PSCb48FwZ
DG+kHQnc5cq62XjciP0p96YAk/cdAuhyIqSpeA90XIXsA8pJ/5OnDhUB/QDZaUWa+CkKfI9F1ApH
z972u8p0Qvb5hBc1Q1p4eHGZ+fsD9TvB1XxzNj7rUbyNEKoisuN6Z/yl91AFSiTIXTAlTBRa/zyr
AgS8Jqx0nMZ1/omTxHPMj+ToVnR+Epi5nT2h0kyWrYOmReRXX+c7ubwuBi0u22jL+ln7D3vC1ldK
dU6pAU5rSU1KXlD70mU8/PbtcERYFXcm9C4h89VM22UnaErSm/fggW76vj6SlLebHE6rM2M7HfkU
YZRm/sq/ILWhCI4uY63ln4PXK+XauoIkyxQ7RSDloxPGh495in6W7bcpOXbQUf+pZ8Jlfz6wnaPq
wSKmbMc6GdhHPJOT9BkZ9Ma1vF7jc0y74tYGhr8hR0ORMo4WQinxMuj07gUx9XXHnS8fChL3LXLw
Q7iLYjQuPbCN7XfZ2cAAFFw2FOXSO7N2810yc6UooVf13DjB2763s8wNKd/+g24u5xGlzxyRbG9A
obvoe0XMC40la1pdRMsIazdzoCDQns8M++wDf1DDE0Y38AdbKzcz1T4023Yv6e1Zc2KoYboTm1zm
s+RQAySmi0vK8E0ab5+zkkdPwlp6oXrc/kiY8znGbA+KiwcxGcSPCiGvqe9SxP7xVIFijr82405l
Gd8NHCm/+jI9ZAC5SGApeHtCAm2YR+h3JRFaI/Unm3oC04ICjGvkHSnQ5YbvvG+sZYpPn7xAfG/w
so+tGkEyqtjtRhqn4KIt6oRwE2QPfnsvaBV8KJaN4lrWccAhyOSwMfmXAIk5oMj2Vky7N8k9Bxv5
6e9E8lGmxgfwtOq7lubh0VgUVjE/3CgmAHK8x7qpqRSb7IanxHSW4E5pZikxkN4WZYrQLONMybct
m9rALRw9SWhzdZOf7zkIio9dDUVpybr8cpOzz7322lNIytFNxixGanNWbw+BHd/u95peZSjoIx8S
p2fXIxZ92TbZgf3pq02/maS9I3BrDdnFW2zurw24zLTn2sdBeZMozcP6rZhqO6LF+9Xeo2klNQAt
hq3OemcA9t/24/msk6hbxRc1u1lDmlEuSP5hNpjCDBy3GO5Yvg30ad14eSUgeOPH02leTuSRNjv7
NwnTfFHcjm7KD0jf/h351/FFz0DriLPNom31M8N7u0+rCinr7LDm5LOecAz8EhdYXNdWTyyQe70A
7IxL7AUtSIIDbi979Yydi1z0xrmixhINXF0zFpe6fWtLa9bCqpVaGgadOogvygdgQ8L99MHqjTDc
0QMTSLdGVGlm3WrTHnugGHz/3AHUIMjcn2qa7Rq07jD1bqYg0jEKS05sjOLBXUa9/Ckf/1abaSx1
QvR0ldqeE9NaprOQdhWRUcf3Px64lT3rYveQW5NHMl9tSCj7xMJ0QqBsVTa9Ldlju6YR/wPcASS3
iROtBebXzMEzMRyL1nVqLFBArSqFzxNkN2Hb6fdTC9ElNm6XacYeV/MBadxLK4i2RlijMbgYAujF
NIaGFTzfJXtj3Zk6aan0oUVHbTiYmPgBLv6CNKb1tGt1m97IQtX9tMcd/dB5jJ7sP1BqBWVJBrHM
cY+rxzn95xIUpa+zWJAlHS68R4E1FDkxMTA5FxXQ3IDTZzfbt/JR2baXP9bYIQNZkJ5dN6GuRu1r
gPMIJLrjU4MHWfHH2vZpl5WNGvW1kBz1TVUvz7q4/lqD/GmxkqWxNDcbFl9lJJysWOEzHbreJWDA
t3zoBOmo0YzXQbo33J3PHfqA8agsxY4DKlLclpS/Sk3ylp46un9dpoB6zBTb1DiOA1EKl2z2UROA
vN0dFMhPmDiY7lvzTCqNvoyQJoCwNzKweLwvtx4ddZc7Es8KaKFtfctgUPhr7qYeFd5Om+XbDOul
sq8bDoIjliJUCjyG+mtR23lsVXXG3TqYOlpjDCqb9amdXtH0kyE3/6lcYm+eDHb5+8O+pAovhapm
RvHzk4OFPLNHgbkq9Jdv8E4hZimtnu5oH0YYMRS9xQR0gYvh2+zZYsThNM1Fg38CDbOXowMAzGtU
dLdHc1C4gF6l4acS9rG5C4nj6qzgljVIR6DbbwUOm/UTcseGJND1S+OYYHXX9pc40hRRoIYvggGF
o6tCDEcM80dnVR68YI2JDKl/zw6A0IExHzrwmLE3ZnJM7D6BflmKXre5iGyBxkYgGbuHGlHzYEOM
U6R+t/2Q4D7r3yanzsF7Hqxtm1rUdtOZs4UKZoQ4wbViBzEluNNYXL2LA8wcdZYGPdxYXMgsUOdR
ChKBouzRdi0/AhdKXH39zgwCUy4JWYpI5hzgbkFjogKIjQ5m4Hhqpl2jcB9LodVSrUZUg7+d1c5p
f7bN75Eqx/AOfP2aKfEsnbnbrBvnDr1Aoi4iW3nrI4WTRT0wb9v6CILEciltzsVvhkjRoeaQBxbv
x7zkK8sI7UiWrM0UwAwArkaYPMBEvvVggYby/aj+2jKDmJuyXNibo5f3P89RfG90NpgLvzgXGyfd
5xXROCWw9b/S8X+VO9OJjpTOBtuuC1Y7JLU3Y3JkPMFvog3P1zBwVLcA82omU92LzK6NBCsc+Kn1
DFeisGIX78ZcpXykzaFb9TX3vGsLQgNlx1DAXUHbiTyjELeQeQIlnAEERL8BNH43u6f/TVk+2gxT
N10WZcXm5LMmj+B0o0YDVS+hSZhUiVqN/Q6woaOI+thzRpXWt1HoJlTtr/8nQn6ufFqXyzf4qwqT
NF0tHnvpYnQomHjqcGoLhH6hZJIKyTCX2qAMww2WfBbSJ0sg26UE+f6yx77scB8eIYuxOTbSXyGB
ZVPKgGPPk5FcHdfF7+RPTLC6sy0obTKuXnYNPYnPv+Pdp9KM7wqQL6u7daH18IVEyeVohRsUHYBf
35WdX/wO5mdib+n+NBAA//AjdazToIELB/3BVp0hWWN7AtC3iMoqf0OCcVC18t/8gExR3yiid+vv
dZD8xS2aE1/ine5C+ho6CWPv728zYeERFB15Nib3qvGt93ZKAYULBnzgDu0sSYaO2POGFX8ToEuw
P3bb2ritPpV7n3nJfsboImg6ciEXnSx9ZDguomiSnfUbOX/xpLoEwmLeSMhCgWXduWGG4/eaO5ZK
O6P/abNfHQUHJpaw5fFBZlYUdxYZcPaZvUQyz1ldlecTkKeu8e4e7ok83N2GdM8WM0WD7zugEFLO
cOSiHMJPtdS7CFH0xIdm76FX/EqwVxHTi2o2Hr9hTVhHhCQ21wmrcIF1zNC27T9d0BHyZdAeml2V
7qURPCn2tRZheLqJGap4k+7F5fX92k0zQ6ysM8p0WZQqXJBJ+gPSL4SXFmstcCoW3QWh0G+rI0MY
/3niTEzDXm/Y7on4d4egyxyHQsTqLkveV/qM+8z/wUKS9/KZ9b5keQfGFBLdPsMAroGEg84vLue/
VKd5CGR40pKP/mvNzfqz5jNAK3KEVgpVxmBKv6w5Pq3/eZe1FnHzSaaKyvwtx5ghUxW8bMC0OZ0z
15T2WuLrTFL0NA728TUugapRIABPSAybMDQjvQxZVm2gNOFctVhKHSlzmIu+j13IPltOtE9qX/e+
TZ2Wfs/AQSaQkQsx7seNMa7ahsuVmZAkRxDz0V3C58lBkw94DX2VICyKseEmnqIecj4YKh2DOH/J
xPMuxQqHqe5/jPZCjbfvoV9ijhlMElUYzT4AP5WuN8cYuTSXWZK9ytPSasY1pu5LxM4i3JOt9Mb9
FkW1a0FDjlNDWL0qC8YbnLTN9MDVHjUih+/69xQXYOuDgiSk4RUjKK3PCYQbzcFAD2ydkwbrffIz
b3cgxj1FEq6GOmU1VUE7gPpPh5O5sPKGLyY0THFHzVEgykBQkFsrh7fcpfTLG56Kk7T68C4A5q5u
t/36l66S76sF9gMv+AIHv0HG1aPSqv8gUoaDNGchYQE79GLj2a4CbOVmupjiWhQkXtu1eIGOYSWz
ZYyYPgZJDGefuYNX9FHQ0nnXucCw/zvdvPHevIErDi0gwtvsfcHM7u3lfwbhJfu5pxZykTnP9Epq
vjC6tRhwO+pYsFA54g6AWOaP/Pe1yKhjVkNxogEWcBsCghn3ras/j6oLf+Kh5I3UeqaRHeaBUF/j
u1ArxHykcAKgCgZI9PAEjo2UxMuvt9FPUladO/c0MJ23rG/WyPll0I1IezLuI5NK6NbvN4HD0Nzl
EldMhMZNkO1bN1GYeUF6duacweNWJdgv6sP+vxun7FH5bKZ7LD3ZArBiZr21o9lR7sYROle+obn+
CMz3Uk9olONV1AA7QzLT/bNA3clkOMVAy0JpgHdcr3puZ3eEBfW/QZf5fcU20EWkErfFRU+to/+n
SwejmjJMh3hOqbtD6iHZd5zuOu3UPljweTs2OAujKiBlvHYLyC28BcO8yibO8Z3KOfFwpbLzutH5
r/gtizEo9FcWL8yqiMFbtYE8MDOkprpKQSl7rMOf/sBwE07MA9B+4dAQbwtgv0EY3M2jXwh9DfcD
0gdneZfHkeATyFibxh2A7reQtCI6iIVrc/e40fS5WO50p8jC33zJ+ylsJtx6vldNqkMXPEp4bRkd
zInzOA/ljb9wJwCf1VdVZ+41BYGJS9mxggPNN9Y5NXLul9PK/rd/aFmnc2ip8/KJCbBbbCvYF+av
sgUSwTg6W4eVwdXwq5a1r85qS3yNijzdlpkogi4TDE95QCbdy8P46aNP05KUBxL36XJ4cDjCFRXl
x7mdt2WKBZt8NqNrAas6ajWEjcfNeTbflQdyGQkMtZD5qu61KVgVPnLshkE2Ou+/yPCAMuQE0leb
jSzhxJ7ja6w09nfjv9GrwCPEpBiHCqq+hTrZ3KT8oDRcUoaPweTkm6my8sWuGw9rvxTqZyiHOCAt
JPkuMAAbpHhq3nk3S4AReKaSthyB78TTzDPBYZXV/e+iorf+fnONLHoOUwXTe0ZzicUWl0CRvhRX
wJOS+7bvK+3hrxnLvIHuPNFYIPsPiu3oGIhJA4tZ5rm0htiNCAEeILcM7bW9rw/fbwlelkZPPyg4
C/YxHhJvq1LQETsZnAIXeWGF6b1Qi9HqLwn/tQQbxpunW9A8pET6+hy7m1jpNUMDxDn+wOFVkykX
P9JrThKkyqb/aeqxSlEkOCNFId7L36rMZ4mB6Jzgj4PbITXO0en0UJvRRENTws2vMlER5lt5HBPl
ev+chZzeMjdBEK4ulL3ndtvUuTYkXFHDEdHe80TXLtjZZzjc/Uii/D70IGwHr4EESS+tkHVmdhmS
sdZe5UgHp4anqxi4B0mPtGlhyFIKXmkAeVT7XcRKDNaG1ePtgglgXT2MXeMJLJ6BfBagwGg3JtW6
rJNCKysmW33A4IfQLnxMuVqYv/RGizePuCRkEOz6e3D3uxz26dZBo0HXjMpsaytGcY3GW1UK35as
9uINnQpAR80qxsFiURpsNGf8ZR5+tuRwn0goCzWUiLTrQSTyucPg53aIZUda0aLNuSTpDah5haSX
puOPeNrp4PDF5ExjAaPvXy7ZRVccFgaACC1LLFwcTKuy47Uk/716OsWSLYEg4aGkA8GmQxwFu/jV
H0qfuZkK5+ErBORsa+HWw4EAsRipL/gmzLgw0Hs0rvJwfz42s5oa2tF6RTAjCPaQjc10JJnSD2FK
btNH5mzv8AbdynePGsnT12iihBX0eUUbQAeM6XhTEhRheuT4467dxZ+0XshvGtGhJ27VEOIb7Coy
8ZnE2Yex7YJaHUkIUzi9aA1XnOsSBSjIEUGteHCgTBm3DzSbqwOZJXtRkPMZd8eS+i/kWnpDwKxx
cPAunnxWPezNOkGgRxEYr2IjgJMGgT3aVmKDTno6YUQ5itCpyq7u9m456FeFvsxfXsbnw0tykLHI
qxXCFwjdGbmf0h6RkeY5tiunxh2GTy/iWdYFQeqX322T/GCgl0nMe48jCKdeKEKNdACfsGizA7aN
aMuDt743tbreQ3FdJkprNmkjCZ3BbDL0L8VxXLfpmBUrl7ZIgCXucXTmd4eLCDYar5m1FdLqZKFu
s1/0QqW6IdENo8I1LCEqSapBUhfS1D8t3VDW716M4dV5OsBfuGhip/OqZUkzq74mVivSYjOe3r8K
pOrBvan+8LyMLOCR93m0iWia5qcUbroKQpBqemOmWOkoiU74O16gI0BsCfSbmSIsxh6GkXSv42Md
1SeU4oT7TEHE9/4gVw6y82ya/z+i/Jw3YZirQEnEZ9GzNbtNwvvEPaRYZpJpSg1yiiAOMpbtyOzl
70YugZI/tLESheQtAqx8QISfteR2KaMejmq5j9gUYL+sc6UVuav4cYzPMK8v4lm37xC64P8CfpP2
sD4+wYB1OaJpkXSLV3/Zmo019tyTJQ8BYg1mBukds+UdqhAxOI3oS1A5QBgeYyUOIULwP4vGl1NU
VGsijqsfFxvyQ/v/4pm4AfvNSZLebFSUFq1XIxus9EsPjGFWIF7nPT8aRxTCuVvoQdsN0qe6xtEF
GACGOPBAUw+txG3ldJ8lKTedZCsZ7D9Ngcr+H9qhnQUkfxqB2ohe++Dj3hkwq2jmFwJtPywVEF8b
oKaWLRiru9TuZzoum12JuQLDR/66GDxOUA7sWq0/ieXi5ALINxaqJ3BxDGw8xnB4Thr+s9Xpt8q1
DvTmMd68wj/sIXaOLrOrPt2+X78OWmTrwEE4hvAXnRK2AC2HOOhMhptogrooH9WdPAfX3sEcxWBu
v+DlmFO1NznyGh26+EHaKDJshn/ksRqM97XtsQpWej0ESDDVYs5Zee70Pu0+I3Ps2CLlhETvTmCb
DNvcIL/dcS2NM/1JPKg0+vpPRxxUjEzh6qbMzFX1f6pQBPcppkHwCeMPJCuBoNN6wuqeQ87/TEVz
PSTI1Y9WWs5SWuOCSy3Wcp7WXXu9vq7+ufNX/WAju6KYNroyczSsUjFYLgouy2NutRF306bRL1G7
1nWg2dEeIeYUHgeNIrbrchSNHQozN72OxQTeuPMAwqvwNIc9OKyXLJZWOYXXSuEr0sQr5hgbglgs
A1BIPJ1Uv7z21R3jsvs2RuUBJJD5cRuKg6eFP2oK+LcggWMi0LXNIE4vcLPQVz5FvizG2yJ9LUml
P0pjHP2IXgvyz9+tdGhsrE2MDDNCVd3GrrGbN84xiu4WqS4DBCBtBy6hXHaf/0stpJ2FUYLi7Quq
WQZ5JpSuMjXMtAH85z+Lu1zr1C11L/7TBEHw+iIpTgCVMUGDNbZcscgWuFM1bt2H4BFO7HtGZS7S
6f59xwXB5Bs1mVBzGyARj7/manxmObRHi6bu3DIrlzIeMbBlChInLst7paz8vZLHTQcq/Utroesr
vO+wwt65k726li2Ev7jjRWnq9oan8JsALVONuLc64Vdj/awfdCfGqWycZqe2lrK2sln6py8TOuOK
/JGYj4pGfOBhHmYTfOLcaFmLrd2GxcrbgxanAK5Aeu04RQKvoFnCfrYQnNFCQ5R1yTYKc+XJJOq8
sZXnn1Uh9MCAHmmhkcT7LYq2zpv7RZ2mUGvTmZ4p6xI+RCIPD++RAh96bzzL50bv3KDwDaD0NXBA
tHaGwahWGlPz6Zl/u3li+e9/icycDYfq+6o1QcOBOd6VhXIQf7lXpau8kMXjT57TdxZ5POCobEzD
uNdXs5JM6JFsCKhw8P038CWUtjDzVVUZslgIohGX6FwR8gn091zP7J20lygxlmQdyu/bDrtN6nTO
FoWGEHrQyM4Vpi12gBruFWYI0Zf9CylO5R8lDC2GL0VsZv8I0rGc11UvLRAs4Ozb40X34NxMGgn+
ZHDDHXL5NH+zA1fZXZ7wCuDzqW2SEswsi6Ty6w4l63kAkzsNKlaZ2m6Gt87r0cBbbtsnKJNmKDAn
y1tp5U22VI0Hq01gJsDmYMBIx4zKA6kLHx2E5h3WkZWwW8ughUnJErv0OQwPL0+gpOXZn7cTS04A
vpYT3pDJWG1lewVsBmEUeI+WmILICnMZYzACV4JRVzsvbTcu9lxoUgtRe43AQPJUZeyptMnzeXMv
kiZajntNQuEZFs/KTGprq7VndFyZ8R2zQgaPjsTHe11hxLKCtb3TzpbjItajLuRi2dfdBvKnBiG7
A43b98ronUMp06PU7BlOV94izcVY9OU0ATZ33/upelvYByuGwp5CnirLSecLuvJ+N2KGKd9jLiPh
XLS/DOVNpAJzLtmSsoV7J8LcWwcl77jbs5YKnZ0tnTYEu4zIN9Oo9pAc4LR0qjYwMxyxx3e7j6TJ
nueEP+GjTOfJ/XB0JgYsTcvHPHOIZyK7vZmZ3PvFMrRs89Ehxee7iQ/csQrXNF574a8lzQ/sA7yR
+cMm9LDuaTSm2Vs8ZhHZ1oSsY5KnqSIVNc6nvwELT9XMYF2xAAbwF42JrF6GB+rZ466wlJ/201iK
c3dAGCfM+YJ/p4RD3Ns/eXSnzrqHCRirShzKPs7FwLLsMfMDHHNDpX24gxo7Evnn2srUmMH+vS1z
ZY22Rmc9pU1R6DDb/Aafd7PGaCrD45qev6mmy22mGLbQgXcl5ZsjxtGsE4GdT6RTiXjaY9PpBVUx
tYZTG3YBYAgct0VCkx9LUzGblldVQXhlVoJQhCAxeMWnB9hpzBVy72WjVTyQeJ1m4Mtbb1N+jRrd
5thdKnFtPKBOgGkR48+a0ztrnj3mIzWNM1O/8UyDaIdNnO5XLbvIXRZPX+ccYp43VyjHU1vKD8KC
6EJvqz4gSdDq0m8NL+15bGNUJKa9E5zTBSiZzVM1ZKnDbPNyNAuTJkxoVvj+3BG/i0Nxe+5+A16w
KXdqPA6lG3Bzrp5DmQMk4kmAqB3W+T+1mehcXx7VmjwZyDcgO9Hzz4chBao1e3xlBGIqcYquVqs0
GGkEivkKA7ATNsD7hmjt31moNfPC+2ajtxzusIlv4v/I8rw/m18BFfdCMHgN1NHP+yukht6hhdQK
v42HkoCPevecp0Rttq5q/SGfFM4QGFp+DhGR7iggPSZVzSsb9QSGXgri82OXG7xVzkttRDEvb7hf
j2cg6OidG8LBh54m9tlTGez7o3quNZNX72Z1o2SqDsahCdVZARQzLdegFsij5z3gGj0mZ4ZRaUNl
14VyKLhta+JBva77ecpqaaoketrf2OiH7ZydidUWBl3ig1KPBNh8vxbK5wzVwrtaLhx+RupjWpeG
uY+jbU7abHgbW/CQMymZqfe4VnkrrJ3q9XW+JiFlCEJ84EgjG5mNiMqEtREZFP4yIYT9Pfa01BOQ
ZRf9dSg+Tn6PONDldJr6QF1TYFJtteHa42fdjlZyxVMZyhbgGYP1keHkP0zTRhsLDaEQxWmTqjla
8eVGJ40SU/Sn/xr+xX7bcH+i8y71DEsAc2BzBd8ViTjPY9mtzZaYi7RVqZRvFcdtk39Fji8DzDXz
dMRU47iJy9A7X/Cnyb4TkV2LYs8q+At5BFDBh5w0iuChzJMGmZTYROi39v+bfIwEGEM8mS4axX35
Ig7TanGadjmbAoPOyTnizOESAtyPtPyLwCt135XKlTOYKgCUXWqFymBlLnvId9R0sL3ONFUxgnFn
kq6v12pl5xkWrp7ErU1Bl3qlapiPVi/90YkNqCKrQUcSn89KORGyFH147C0wwO9dH9mYQGVRH14d
n+MYITpaPrc5zQ1GoeJBbowTXk50FTfAfueBfMQFh74gJWcjcP0GfQEgPAw0EV9vRgz93eiZTMbi
JNNrTbZdzB6Ovzz4II83+g7VDr5MVu6RhkG7wTovTB15BwPsAAi3xRgpGcLB3ZvUEOeSdxYNgfqr
w4/18hVmUaP/H/Owlal9oFhXOGE/bZ8mg2oZ/8TKMsT7HS67qQX0pkVo5VAIOJW8mMAeyGouiqZs
Bv1LVaFgcNwRbRHKawdpmUnvXgBrbpkjnw4V8jaT1DtD2GjGwdNOWooVZvNw+Zjj71/EopQmgSN7
wnOMLuuvDDJmRp4fv4pVFd9UPOnUQoJ6ufR9OJsUglxKl79FisTAYxRdtZ9bxlZxpBlLHSF5LOz2
xiZpsddTbuq5ooNRvug18kKlCRO8NKItmugru7pF3OKDn1qu239SLa0KkwWHopOPRKV/CTGIeF4Z
LmA0Dt8bG/GqciqF/lXw+9dWDssoLnuv41oAjynAA1Vm/ZRA8kSr3zQEqwuHTCoSqEBEFH3VEqId
bIZidG5dUxB1aXuFvQfA4Ucf7UZK8KAYCXcdl5wCox6yrP8zK4ebjquw/hBSHRvWt/y7WNx8RSPq
+zPU1eUyhsoY0tHEzotIM8lAA0HTMYOfhghYAwk7SOnmukqCqbkXwR9YmbfZ26+7vPIoF0lwTlRN
MR+Z3ist4Px4VpBjBERP8L0NbhrfsQO1Z+2zULT3aX77AOQGlKZTK3POuu0lgcOLetzM38nCePTv
92kwvWnQOgk6f+mHevDswxSPvLa1YVcGO3zAKbtqayuhEtSenz81tHEsAWMFDdFQEYQ30xzzuwQH
aHgdst1AYGU3lgUIsHL12wUeeY1JPWSSHi4KShNkUw0YbnAAOTnt6llO5nrq8FEljCZ9kH6UfjVu
mbBkUeQ2Ddttm6yqtpOpJdQByxO/ZzNxW/LGSlTfWL+MfXDJFC4M3kjujCTrv3aYV+xkrqp5UEBH
0WQ2ODLC2RfQJP4VgfdouDbCc1G06Iw6jZStNdRudmmIKC6X8RQdYVxVIVJbT79Pf+Qc3VUmw5zb
DY7JFN2+PyUfUpQzYVToyZaweCGMVeF2fR5fbRH4lnUHNdSYEge5KjP+rLjCPmz0tocA/KpBONfW
tTGK/5S+Qfq+F9BexjT1adYn5dTQzmW2MiKZAEPnKLu0rYL/5KzKaWzvvC2SapdgWhW2m5jZVIhM
zGaEVxjb5+D+Qh8EJT3b7AvytHf8IlmbQG2cYOWGxdyEIPI86TcWZ+LN2uNO9jE2sE67Wl3gLYnp
yo/7vIolyFHOmYqoputTQ+1y4ufdLy9Qp/svElFCEwlCcZWe/FTt9uZpvDHRzqq0FNquTACEWkNs
PcD1hxY+ajsiYebnRtg4E8n9eIqepZIUIvAejldwWFQvfIQ77crNBUXvJH0VUjRQ+mo94+uqBafW
rHzvfvCsErbJbkcxJDieHF+/EXZ0rRNJd29kmxbdeKW79AhuseCkappN8LFnqfM7kRlsBresj9av
GTiCkt4KZbCdu29OLOwmOacTUNxzfmUMBGT839BT4Rky4NCMcbov4USL/s1MRQGl1zHxg4Vs9Jt9
xrNsEHlBc8dGn+pAoOZrJaaXxorewFox0s8wej3GjuPmozLJolfgBQd/vs2nDU8RF+BP//qLyCce
L3P8cjf3cLDaJk2jyu++SQco1xphRlUFPvgFDqxfealdn+RiUS58DtiG8dpI6EipsXs48pWT3N74
lqdTACqzZPvXZUpMOIbrKcqKL6NFLy///epOnGX15eiz7yTw4Zp7Cvnp5IkVWIxTJ5TEs4R/WDLt
La4opBlV5202wyy4X76lMo5iI1NZQJ9AjTEGHjwNXXLPcDK4hD0lPPa88o5L/YHhH5gKtvrq5dLg
QZd/RvgAlzoTOP0dPvnKc10vbGidm0em42CHU4J2lE5d/ePnvbiw/mC88r0P+oLQh9DS43CRCXiy
DxrJufO2oqYL6PR65wPeWY1H0Jo7TAOufRhH8o8hyq/6H6lbBX60QTlCFGG0dSMFORHvsMJMsjU9
HNu2wtXawgOvxWjS71v6Vs6SlkbYWRibhc1ZSKxgYgpYs/jcnCwwDSx8TbnUU5IW+G6LR1+QX3Kt
X7nfBH6P7+z0YLNdHOuefvmf0K+N4qBKLzTCriwAbtsryW5Azz2qKWhsw65dsu3AjG0ht7qmV4eN
yZrpfA3VTW+bI2T3i374Idrxz28L47GgxhfL9viNU6tdphBXkagMmVvqJOl56+uhMdJl/7y+Ymd5
Z03+FtKkFFJ6SO6KohTHx8Hh1LrfrmOQNTm/jmupNogmIji3cDfnbYqtqttmkxc43zTfTyoto5dQ
fXRpEOsI0zb5rB1ZdQR7m9dZk58KdECYEXdwM8xZSEvc7q2xh1jgmGWE63OjJkbStQk0g6o8V+EV
3cO/nvL9HrBVSvjuf0bwjAXuLSDTZQynr2b1cppr6yTBNd7PnocM7r8HcNYu6xPjFd7L9eFzYbG/
BF+oa3BpJVNBGw/PEyTEuQJVvtqZA3B8iZx3vgiMQ+gy/2FnlglS3wyBI9oog+JMSbwXVZfwqUId
/HfmT33m1nnYu9CZk52V5PwtZxpsXUhClKNmJK9Msa8aEMiuhQaaNvsliyY1yuGPYA8FD1cGjxoB
m6uwRcgEfUMMxFcEEJVUVMmmWXDq0X5/JVP6I/cp9Cjwae7a+keJYSG96Bky8j0KxA4WyMX+qFDw
wA5KjDMLDxEd3qmSnxw1KzfIgrGs3W9TJPiKC3HCDqvy3lgaMxPZwTk+psZViwQgLGr3c4dLidYl
Oq4TGmLHUgL/tWFLhKDKuE6IseY7A1D4XWsYNcrnfU5W1EIwiScQEhk1uCPywxK/7PErYwALVuwI
oE0TnmlfDPnPHkclhVwE4ojeS4hUia5zLCmfL7TqxWw6dANb9jk3LcJk8/GDLf79/dns73pxr4Xu
h7uo47WTepnVBJaJ4hJqqhPBgrRX1Hcr5Ldr8ABETgpoTkvVrQTtCO/7uNV+f+OlhdFGnGp/HMxX
SHNDm0H9BBXhpJLF/BCULb7jnPj9o5q8xy0aJp5vlklDVZUXf64c4cKo+M49YpQdH4zCgCNrg4fw
7Ab1ymw0ptH+qK1JPWstjvHKs9JIoje9id1+CEDNAndBncJGHpEQpARXATWIR22YpsXB6+B/XtCV
3E2GVispVY8/yRgKu0HdnB6U6dRPT0j/jwpIeBa965kako6IKs0Q7pKJwImsjAKSgwynM3izgr3c
6ngCAivBgGIp/eyRBDlTMHdnl8JZiLSm5aUhDztRRXXz5udnY4W+AZQFcVGCE/eWVC0bgJpxc9NP
K5LJOLspZhD74KW8BmU4GWW+Qap3boOZa5Yu9pD2sreqS7ZyvkIj0SsgEw0WqTrqqVtutTRGpeAG
oFG6na7gBtiWo0rW9vyEe/MVYEicKrKyKEUonUFuCJiH5JwnTRnU3ungPU62z0towJFiXivgysaQ
+xasp3i3emCMA5ME2+Eyup/Ad9sHtdId4VEP8seYgAJStZyrZUmnKxtjnPJZHKV8W+SqBD5+0nsq
btc+QvCYYkyLi4/tuLfKaspN0vskqVu0+UnPm870RMnYMtZb++ihkwe8tuM9on6Rr18EkZxJobFd
U6GXuLCjuewIbdv0Pdz3lCSV/R14FCenH41qiQVXMMHO9dXvtokz32mV0ULcRWyI19H3Fw8bGTVX
6Qh6oGABF4nJSNW+bPgXx9BqD1C/Nw6ZsnAoC9IV7NIMlpAC5+0VwBHn5S1OiLGWb7/5Wg+wSmTw
oCf4E5bDYzgfn9kMsBkEpkrev1+eoAVRJaw1VgDtQbcWFqvdSvbLyGKGz8vfx8EqQTWa0rwmeykU
BO6NU9Hl3ySngg3FkttVXkcnPsGvX6jAQSmxNTq4W/DCDEWCaUrXV9WtAfTwBaglSG54BTkMUkZO
X07v/VjKjzD5uz03fOZ/+nI2Ks0+1l8T8fLApSwnfvx3qAPOWMuwaouOX22a28Q0q+ZbG1tqzAdv
MvCr2Dt3BXfuoYCL4P6z9o9MLqnndNwZKdtRqy1ZenyWhhgdDEsI3jzUttI13zK6K8ZWKB1B4y1c
idyFaXomIlxd96Mth86J1hgTaxDClDBTDfaXVV6jgZuWmkr43ndi3SLEQOnulzvAjKspCx1TO+3k
jI5CvGboz+GGN5Q1foi/9zaINHfFWVThnWy+4Az+pC+njYpp5PYyHjQKySCAbPhWvvYtN7hxNlFh
xbNVbGgn/Z/WFUFuoZNOZJ8UBPDQL7gGWv5Kt2Pq9FVI15D0Vrt8ctJUiZkM4JN6PrGeRVtAMIKo
xjEdNQO3/Izh+KnqDaa4Q45WFHYnc7omLYxN9uFWKiJxEul5KIPqxwd1Q6uwE/nq18uXYm+6axXW
HXpxFvj6XGRn2K69i4Ix3XamPaWt8tVM3d/FyIHSPol6rBUtRkXO/ExBT1Ww/F+ZLLzRYoIAiuWA
UJ17QCFRqxUtYjgvaSpG3fspNbif7+OBJrF+tByuPx3HCmdTBVCiHnCwi6y6gp9DVrP18ighjyxI
Zgj4mbqcXNRMmwzb8Fnm/HYAnGUP1PMVmVGONpnCxAj14p47QnNBkG3xZNXdhw7YO7HP9jBtIJTh
XMmrsIhUwA7ljhf/cQ+LhZ0OqFvAC8xgfwzBXVoNg4nlCIwcYUBieH0/SaFHjeooZ4ynBnGo1ShQ
63VTciHQpHadwsa41IZoTZSR9BC3Vbw2euDAn1bDRQHjYWymRsM9BC+5Mas8vyrqPPL8TmX3xV13
OxNZWzIflijn5ysLYGIooiClM84ua10IqHAkLFAesjbP/M9/h4ttzrZDUlJxAnc3mH8yIYX2NM58
VdX7yWBjYEnWigNPxGKNiieZVa7rs02wsTr8CzBijlQCFW5hxAinBMVUi33k1Vx3z5fQr6s9hhyF
4TGO4Rh3j7DQzujGGOjbbmXAp4xUBUuvT1ULrVn58NQsZQz3Hq5MCnBPZm0VN3Gf8JnJpMhiwN25
qRXX6qWkm9Btc5KwUnvRKGKIrysOEQNpnehrhhoxZ/JXis0kMhQBnqbwXzKVgTvr8MgGSvI5YiPB
PxeWa0M2PAHZQilSAUKtcjsdrrH+PXn7zjdSaVKoWjB6BopY43JndCyuuMtbVykBGaNYtjdK3tA2
/7D+TvmAup11yRWqn0dJsebX7y071eSTN3MDaY+yH9RixTDIhSGYsbK0p20YscXXRa/LJQ1n1deR
JhHU2zMOA7Vgrb9O496LjXyhlSqYvWPxKAD3MDLzsmsS/1W+g8b0yZfDNTkmcqEbMNQJwLpd4ErF
4QRnJ2o0kRihdiNyOM9qIwlNRhSLu4iYVhYGUhZ4BeIcz4kQtd5DYsSTG0JgsuXHOOK/px8dXJe+
6t5YuXJc95BnSYrFoUDQP4ahmvPyYIpzYvdwvtinGCOBVEOaRCMtbIt0L80jhDqE3PlQqw9p55Wy
RH6sacFXnoAzalDYoOdXQlOkUhK2F0ueqXFLrg98eQeqTm8XvSKMiHJzpKi0VO+MVveQl1ZM6Nqy
ySt0Pz0rSfkAccEezfjXLfSa6G/ODADjiconreYY8qCELEENP3B6oZzoAHOq6UdTux9ANB/cd0+U
QCJ4YsCzR2DosZZAOv/Mdt4n/6zZdnv1SWSgja0yx+vOM/wbUjCmC0Nv7Y7JCGoZJzm7HnxjP1bW
hE8T0XB5OPYOh7nej6qhKcfsr6DQs5PTz5u6ep7vTfLPKGQiy3odngwDb3TbEaR5LnehjIS463ux
CZSXas3Vm+vwYQ61f/ySnARQ7oqiUsHPn/3/sVDQsJOW17tB2ZucUNaHnb2JQN+nF+0M0aa905RE
2EMXDW3SNzxtWbHkRHeSzEToelIiF6Ooe6iX9bYrBDiCpDJuGotd13SlMsaCZPN9GHNPSx6qFv8p
9ubcmuESM4hDQwfkJCU/tCN/hQoTBC5+wIUB53/MluwcKuU6LHay+zz5udPN9m49EPOuuDNJa86+
SFFBBr9nU34/1KBkvyKIHwvCWgwtElONoa4C093o383wRb78m8wQ8W7ULMmxrtDXeTdTMQ0+TV6H
p3c6uTrZwr61MtWkbvGmCFa9bG1whxz8s7v2w0YwJ3smtfNG+X5l6CpoenMQroxdUdpytUaLXsEl
VocT33Fpt4+qJoWAQxOsKsFw64fmbf7pXPu8m1i6KqbZso+qCIQlZdJrHiOpiQ4+CY0R1CnbYc0H
+jlFyYZ/IVGTRdMuDtHedadIcpXbSOipPs0vaP4FPv0XEF//7Ta9zcndanTBLp/Q4o2Es2Z/2H2S
8K0C3Agz9GWv7jRTPLRi/Jqa/g3oRqJmFIb3tSBSz69kTvaxpmtdc75pJNIdjAklBoZoZV8iQTlf
DMSYhK2HwhIVwurT9BMuqmjJtWqLsiwOY/kuE/6rHT31Ry4CyHRsuqr0WDfPF56S/TQBAIi42aKu
vbR30nPgVYPug3PnQY3AcVoJQwLBzy7xzf1f5+lEQB8yjIw2AFjrR4POKC7mAOuITAF73FN4qNLY
TfK63iB5lRODPJP/bMQyhbq51NPu/874Zt7YFNbRqJ8AoG/heq/vrVp+z1jCBUCPGEWE2+N4TAOG
OuT3oonVCFj2EPgBWvD7s/V004QVx82Mc0QiTBRt62kopS3fCRmEvqyYO5d37VXK5arPYGBCdsx1
jndbHkDp5sxpAw86AbzLYiooJaYbdWIAftGl+KGNvMYxr89XsZVwP0ZCnPzk4wWA5s1mxRTSvqoD
piHVKbbeuS0T7/U1Lik7skdmQWPqcP+pbqXH2UcmLQS9TthelAy+Y3HFdgw7GFn46MQ6Y5Nw8ADd
EaC7e7pUMrNi7aLkL4/HTIAC8vNEL52L5QYmSezgkQdb9hOCWHsyZL4MIDQcUjyfJZocMPSq+LZC
t0bEzc7jE1WES9dUS82fkPdV781jWt9e5grujRVA+DCSwfRGgntTeuWar5XfO06JuP3RcO8fP7Or
tHynqYoE86mjls9VkFbfNPcbI+UVQgYkWnk269Clsz4cgyJDytDonzOQBmUS+NLk4iCPLRtnVvOb
SP0mlSUCNfV2MZ6tNQ8wLe3TjZNTWl/FcaxmikTQ0do3To9OghsNkz0xvubaUTj8JrxmRzJdXUaz
0Z6Bgm0eHHeYxYs6Oub36ZPhibZeQzJiR12x5s5LWwYhEFf3FdizQ/tR3u13LgjcXkuZq1d2leFW
G3Q7MlLO5s1RdFrOBm6Js1wuwVicjFV+6Oo+MLHAvIfJEg37gyRvGkEJAmEdw7qVd7wP61Ss9cHz
Lmal2uwI6ecmmknTnBtQsRrD2K3CIKUAJftpPfZ3g5rQnzmkeUQTV9sUq3HfsVLh6DNBiutBH2li
nOblSZPNh8pw1gs951OUduxqLvnwV1B3wcUxvsSLqwIV/hpIG0Smt3hvr/N9GDmxNF78gYAQpWvm
8H+DZQSuPAzZFyNfHAM/I8WlQ4619sFb7GFJ9oIfm498WHIPqUYtasBMyTraSki1R1guk9W2g8t+
Rq+7dMjaCNzSojhS7gddz2lO/lVuTMa5rHkxCBmTSJIewUnMZ9I6F6i8Dnv5dwKx7Ld42OegSkGB
j+qcWP2NubJs/QoTGT+DIhtRiM3FMVzwOpAge2ZNrl8mmR/biNcwq01sTygmkSVlKXzq4eX+uPkU
O2+7UW5tOgNkxBCNf27sZPGrFzVOW8tbYt7UDWY8oW6N8mRjJiTXWlRo8lebHvKy8tzLI3ju4Bec
KbBQK931DfAHMK5iMmDJOd6UoN7qV+jL9CDFpEdlRc3ihR01JOqywJYfaM4bYlsLXZy+Xiw+fdqP
0sBp0o6kuy70zlR8jwTdqrGpTm84AelrvdQXsulfoTddXi8+MOS2/IvwFFqKzyZ5+Dg2W4linCWx
N/MAp33v8CIAOqfxhjojbagsJ2dZTuIWTMFOvq2nL60MhZtsPpG/HUXBDAEOcYkeZhp5UAlL4k/Y
2NUc5NCyy5BRuaTzGERV9Z25fo64HZ3WdTJNkOmXBi178tjr2dIekmzEJk4ezI7IednGr856atDU
Y69fnel1YdRRgkwDpsV17qpQvhHGFcrmwMCgoN5EbTU80pWaJdpnMBN2fusXsPrDQIrK7gHZVkBX
Z1DRvIlVSyNsNIPa+v9+fhC4gvFWg/CETHgiyBUsZKf/9q59BXlQLhcEi1ttKUWkUMaaXWiKjLhJ
k4unlcIo3KceRb1vFX0DBSawd7X4gcEwTnkmYdeLKHPqftqgtgtYdAau7/l96DkIkYfC470D/vxR
iW1epq8N7u028mn5ZPpvZz90w3Pd6NRnyIYnK/Zt1BzTTlewWeXmancVVQhcOz3nna1SnXLzz5Gd
+YuTNg+Ypxl8zqQN2MP/mQM0rlAwcJmzFPRo72rEMkBGA0tFbaB7KkMwkxH+E7wYlYh+wdaOdMbW
HV0XvjhNolZbxQAyVoQyVXFA/lKiZHqtz8MQBqMe+HKMHrf+H1NpXKZg+W/J3fkI53wB5vH53xW6
uNdGwemtcU/NKGH1QNNa6dcIHTtnBJPCaPpEZvAJhgPPOwA9Mc4/mwx9tfCD2HkqqLb7uRV9eum0
Aqg22x5lzUfiUrIbw7+fmeGSacTF/FQqRiZJq6GApM5sgVvpkGWxQRSe9XlUSFj1oLx64uWmnUVX
h7H7EF4HIRwFsDMoeU0aK+4x4xQfGHLhpafRSxx3WREsPMi4FpL/Rs3yOfblHnAof1NdOd4TU5dp
/1hZfavXBzEMvSYhFtMXG3Spfq0R9TGuDmssd8frMJpBEj/fUWC2l6xut7PFHhbnVEwBXFwiljxx
vFjQYkXLlfuADKEGKNgLlbJEgsVxeq4gOej6sGDAobHUDIfy/b3YVjkTjainzBDv++iwbW2jLnMg
9QkDVX+CvJGKkT491z0h50BgYeFiVxyeW4UEVqQIMBnhubmGWNy7bDVEGZpPxJzgVDyudIhp+xQm
jCJX6sJhiHqOkO2S0q5RDhoo2XY9W0oln6KnbbM46uXIlpDAe/j4JNayNpHLHnS1Mib/wX2a23Vf
1xSLXDdOojnaIns58571Jstt0Ib2CRm1iBx13eqQ9/sktNXuGiZ2Y9e87RyWocSblFwVnTh3CeBm
zeVAatBfyz2r2mYlUmRJeEltcIdknO2kL18CirtUdv6HI8ibpT+uLuKChKhRfyimkVxwAbazWSX+
yrMN+opf3Y6U/xyVipymejhmK5yA3D75a4Fvg90E9MCVMVWW8qT4zmgoJ/tIFgcVbIg3bBTr4pcZ
Wr6LGs25slcsCn7h8h/H8v2Qv/nPnw0j13pKhggHMAOr11nxWGL30E0T2zQ8pvBpiWtsVGfy/z2E
HB9tFoM4/1bDTyfBaV62wQrAZ+d0uUH7h9NALzOw2shQp8k48SqqNWzpL717zwsHmwwiYeLG3Mtv
LAcHQ/F4It97Ap68+3iwerlqur9pSKA8NWWA956rjQLRlckaDWc0fFqUfhAK1lEc4aM7zyNWqhi5
KI5/7aD91olRIVvFlfqObmpm3k6eXrjjkPZQgASncUDNSpHuNMhlxWJvfY8t2VKVuAHcm7A91k1V
aV6r0wjb3Ijzx7kV+8BnIvQKwMDn0p03JKPJ+X/rnHhDVhKjJwq5PfzOTpLBrN7ckEq+kRd+bw+I
efKhS95hSAo52Zu5lD389Mfl0bhRIiQzoYlAF5oLZkUEOOPP6U7alhKyWHtkQpLw4ul3iVS9qXRL
QuXh49WG2/yWRcMg4mInWeNOuvrtznxMZNKS1cDd4T3q7tqLvY8wMonSxNz55o0aQnKlTxGSxiE4
Svz9OQpnJaomdkuf/I1pQ9jdUS7XUBCqQ+5s2+pkZ3/oOCK5on0ONHYMtqA72hKlXHnVf7HZXEq5
myGqOVrzrn5do5yNEWfVCrevgk10me3+TO90qrVvPQA/HZfMN2SIFEb4fWMui0aTdYjvIfkFJ389
6JQceko2jMNQV8ZhCDfLO0xhjW4nZs+gmCK1+kP7eC2H3uFQ6mXjEr4O4yORj4SFtq9Q5mtWLU3i
q9x+0SRLcuSECPZWTRm9EgS7ICfSO11EwOoddUX2RUk4vb0KXpUHBvPSMzAbFi/fCHKqutgX/Szi
0VKtqpRZyqPPiztb758kYd8EJrByCa8FqT5Uz3OE121AXtU0umb7L0omMi404TSOxgf8Ww4iil7j
UIihbMlhvcJBVxa5FUuQM6Qjmq/j6HNlpdllX+6jP/Ik8tbu7TbeYG3eohlBT3ifdNDRoS/nKMSM
+OtywdMNZcld92xKE2KM7d4OJUuvgOOkZXkbrT8QZeRnxvW1uWK53qDFhyC8Vlh7j9jnyice+9yi
qN99lgCkTbtCBVyImq2VjJMVPPo1DPbOroVzYtvAiNiUUWRO0Wz9Nc2CYSPhpyfqBK34TFr+1oQ0
Ky9+++zoit8BvJ6SE0NZM6S27dercMg91J0q7hsv3Go+SmIpy/PsToICcqHt/vROFab9gRYSxjZY
Oxa0obCjPtb5WlcknxuV9EhvDyITtQslJZ5UO5LC8jK5aBTv0kGsDjDW1z/UrXN/3sYYJDHcWcbY
ryfqOlZUufmmH1y2dXJX1CSYSA9b5Q2apvs0r/8Dt1OwOdbHa29wOuSIgJU+pghn1M+Rk91xe+BU
y7WsFkc0vqmcTb0eTsdsukLJMPFGIWCeXoWhXln29sK0VViO6uRqo8M1RPvKVnuEcWlDVutHmqNV
KvuzkSm5RRAxzxlvzdaY3nXv/UXu056RO0r+/VEqILK+y3OP1831K2mV82ZIXR9P4P/jgkvQGvDQ
JV6zsp04GW0y+M3rBwkCcyVSfQIX8HlmHUu6PEQQ7P/AAeCW+1cubUwgpr2CsSivXmgIJseNj/ij
2uoLh30u1mfFMAc8zIxZpHsEQs9M5HFThMq1Ct16mh347so2HKfu7wiEXvBSBIkHHDaCpOTavtGO
lHwW735IaT0uRiXxDBb1MnH0rWgpzJUSuyY6yaz5iFwTgBbiSxQIwps0hwmPslBvWubCmhMOk5DX
WwlHeb65B6NKlhlCjrtMDQ7wcdgqHab2pphQlUHvTOuDo5+X2o/M58ZKGM7Lag7I/wuLGZmYy+Fv
w3DY+DS5o3JZRDsaVlb9wcGPt4+dgmgxJXrHfStFMBcrx43SJYcTduLwN7GZeLdePC2LeezcOs/7
Hqnxui1hfAd8Ss5Qx7tcTOmeryINSpbj5UJvIJQyr9LqZiOGQ5hd+d5r4/P7sz/KUGfXBm5bHRZn
1h7YUvsFR98L1fPFLNGybstV6+qZR2Se3ISYxZof/0Gz99/KwpBYA66KnvYvGZxCUCwyHGVBCEI/
T9mnF5BdnZbgZw/hAYTahRL8ymYH1OIshEqCM7If8i153VhHlMhROe8NKSDDXY4CZE6wTW8/wwm2
/l6MwwvX2YgqRTFWlT2ax0wTQzFaBKGyd4DyxR2W+4TpBEhUpVtftNOgzOnl3WcJxrnEJXqZgQCf
Xnj9eXrOalgUxO0tFIC8gTfIkcsyisp3k4Kfdh5sOMERKFFFr2qvkzYrfXggbS7qhSKHwHrwPy+M
9ltXYcvaVlPI/brkFK+Wz/YFdcPlv8SjE6qlidtayM41ElU2tXmBj1oXYu1Y6Hg9i0UHFE/AR7u8
B9VFmPPaDtzwOxbzkJE/9UkBpR7p0SAbUiK3KEMkfiL7t2D7q54PwgIFnjQafjiu8oW/HtsHwgM/
P60aAEmH7uY4Owj5JePiD1gJdPgOb56Dq0Zr6Pf7ETpQwWw6nica7PxedkTV/9lpq6VIOyCZJuNn
56m7avtCMZj9rwYxYuVF+uyJ9qms3YikH1FLpfM6ffi0QaBoPHWGtNlX/8xoYclP2sUJuFbY3MDa
EAnnOC2TDNHMEuJaE+Ak/EQSIHYuXxv7p0MPotsLIEo7NBURYZWUSdjwRVVc8+DCt0+Owd8IO9CT
8XZzKtLNv6PjV+LXB7K45vc8UqgMnCr/61fX+OOW3hPrc+HB+K7tSydRfYEUAxhZ42PyzWSc2giS
BQoY6zwP8Gm/5ueaFaxV7U2PpgLIMeG9Ib6HhirPLn/yNE16Fj31xIWtCTn0oqFDXbExkxfkx8lq
IpepEP2L3m6nxmfF+3cMesZuQawWgpTsSNl1vhGzTiI3foMXEYPLfSnn2QfA5vCNSY12yIRfmTqY
TxKUNCkId8dOCcpKYjIdi0OtcNYEpwI0tc0CAT8SuLBV1opI2FNSXg0AtlXKn/+32qcClXg7d6ND
A7LqN6banbYeBabKH2rfvQvuD217/ROx25hE2c7ZVXxmP6xFC29hx0p2Y5oYbu06dHpGd4jnWfqK
2Ng8nf31p0H/TK265pXXVS0RNnY3rACLODDsKACyiKOk+KrNUUrXk/NLoriyQCPCmXht506V34wC
tilCdXFJ/zrvfDoPd+ymJEkq9jjXA2UrHEDkBvSzxre3k9/Kb+63qSqJV/rNUz8Id8ZexvFfStHM
hXANyDeBfBUy8gRWVQf91ovXLzDql6hkXi//r7276Bczx0Ck/Tt3ujjHlFO9o/pNxm1nRpj3iFX/
Z1oEyqsx4ChrQSTwu1eFWOZWxEVrn1reiLlsnObpfKUFDeE9PUgv0mMe+IMpKYTewoWJY35EWGT4
Wr9OELYYeQNtEu1DE/j4cUweN9ONU/5eBmWBIHRJYHvW3jD9+iLxCwllhIK/ZKqxpqK6Yiuzux2p
TwUge48hUSPJJ67IVGhvm5xJOOSMEjXO3iJy94kA2gS9MClURzl5i/FpRI0rLtiVVTAltB6/GSAQ
qoCyNEb0+GeLKCEgl7tHu2OmrNM0A+QiCI4LDnhvoKeLfxa3b/rk0atcf4aJvAcdeHKkWxCk9zQC
x9nMPvQFhGUSSRnM23FZLG8SAE1YBgXWGrn/0PKT3PuVze4lTN45ogMrh2OIlPFNDmH/OtlgzSjV
RjbFpU2Eg3xe2uyXu8HGu2cUricH/NdJPO49qKYMm/4DxKivvfkNDUepGSBvOcsqj1Jj4qV5ntOm
PFSI9sg5+b7/JO9mfGQmvvswTr5GASJA8q/s4ZDxLfVYADnsGmBkOsLn2W29enXSAwYkHi13b+5Y
Cg0AlT3fGVHzv+uygAGtl50d4q8tuDEoimTCHe+rJx6z7TUbSHbD98/OPEkkd0f5CM1H2jBEWTVi
NZDYCymmLvJngn6YK/tWKUiwKPWgxmewgfJwbH5uAqTWrbcW9ZGK1v+cjUYdHVq2WNnP3RgBrxo2
PDqbu2G0FbKDYctshlHZ5j8nZ2w1heltzgfIQ8BEzKe55YQ2iYdD8vrs0mMOKgcEsw1/6j/6BXOA
d3NLokR7Ff+nplVEfcLg0aiNsFiphkkF+24EoBgDstBJVc7uSgUqzSUckk/hzU4xGR49x/L6oIN1
vPqzTq+ceR+rvXI+BV67iEwhXN0H+n4ygS373aWSJPuTaOf+C2wxERQaNiVjC30drm8XO4Lu/Qkq
lQRLppqwCi6K21cz9jAMY9IfuBne1UFtOjOi36hbsD6Fl9dif1vbQm9f8rNSmJkTv7gUAovQfqZt
4+1EkYslttcXeJ9C3MXR1hw1t4ECVeNqvKJ0l7dGfGAiShl08iqkoOmC5BFi814kJkxOcGHiWxoU
5gOnlkySi34s3M59rsyFFjjpFKBsk5uLVroRdFrjk9bPO6upR9wbWcqZ6AdnwNOdNO9+r7Murm86
lRACJqFY9bf15Y52zXW7gpgSYUQK9X2rwAbrY5zUsVzrkaEq+LmyGAJZtYbudflsxGxrIsYhqoTp
vV4iJ6FvkwAogd752PnzQpcZEEvr26ZCPLWalrMUfThvJ7VDPRJk/sg9imekPPIkMNA42uoQJkGh
0XscU5/1AVt0hnf8VIX+JF2Q6zQJheXa2VtSTwOiof1EStNXYkglC+Wj8uiQgW+v8oU5RuoYEc+o
IaCVSjvunS6COay9FPC2/RKFVEl8NZUXcRoaJT2OEg54t3RsH2rNS1T8tOwyaqVGTIizbQSfiz7H
cGdwy+oJAiAJbV8qtHoz60WeH4kvvpkZ4XKH0G7rewgxjzVR/LFKFcF4DGRTIE8dsbRGkltz7Hnh
T+yUPOs4J23t9F4aS7VL8mXqPMuBoFUzjy72k1Uwf4ya0NMtpHHN6uR7XSpx66I0DzApnC9EEydS
P3QGUZtSFARbHIwsU8Mp5Gpoaj2jkFnytJ2L+hDCjm9C/URDE52/aERIj+JyVjt7QBTKdMYWNEBi
O9aGdi9Xtx4upUUc77qKaLAOyeD0MeuvPfeBZsoNlYo9DY/eee7v+iaqEQAgvS+dof4hHmWdgWGz
AOXQaYThELt23d3HQ/2B56gTdzqd5qoFzlv7OXlNARBGjqCqeZF2hIflWA+ym8XH+xgxMRiBSUSc
WjNIHoJAEoPuhVO10DwjGftpbEATkHKxRtnIXV5eku6KLz1O2MP4NjDCfPWj4YicH7YaZJCrZErV
HgFOS524Fbb6PAQVqOM3sXoXJs7nDHTnqrITQIs6DuHVIsoLyMimNjfAOER4/CApLrZdI1ZWR25I
JvBQKtkxALwbqY40TO46bxA/sn5N/C/0TP6PJbBocdawilgewbLPfgNlQn4EAnacm8Fbg+1Cc4Zc
6yQ9Vn8vqEfV1LAqeGT9vovm+LPDQzsbQPlTWct6d0Nps1O2XJ4wR2B2Qqk3/W23QZOmYQ+jMWLP
FmhBHB7xhg7mGMLiAQusKsDnGXqci18ygWyKfJSPUnO7lV6By4iyBKQTwIKKxtuuXYnwRJuPLoFs
BXk6auvQtFtF5r17tZ7CLIkRbExen86dS6Z64RHwJwFClsIwa8ZEYHmMfgSGv8FuGwKwcOYIwZnn
xNGQ26/WemvJ10xdUWd/l148zKaK0N0hRJQTOhf7OkRRFkvLw6Hi0zHwrM9tZYO8WBhlXtk9h5be
fQSw87/EJBPLGq+vDe4ANoHmpX/I741z3dHRYCpeHqNLdJAGdfVSMx6C+1BvqZVCwiM7+284al68
ngWqn6rlQOFuaDrdE0ihwr5yPFtN6wI55PWtUvAACELKxypl5Cad3HGW0OVP6YZkfrM+o40PCYid
paRaGg3JRQu510/sxC6Z6p2MhO1Ieb/MVjl6Q05h8BCPEEkDZ1cyQ2krB+44B/JNy7dO0d2D7R6l
iinm7PgjnuznZ9LHI6cFm5j1TK31Hw3z0VDqx1gZ3cLRCFp5IhF5QjxoJ7tjxB44cFWTIOS26wlk
3LBAarWDrKzMoXuCt9DyzcW8qhuwofdSpdwGywYTIOdiZVpYW5k88cSgt8zEpyItCVd5OGa7Wz51
QzH62gFu130Q6IeEgzx/TFSBVz1obNPgrjBKGk05ooY8spmMgUVfkaCSOZvC9Y5TyFcpvMVEYbLD
DeoEOr1gkROdH/LQ4VFSti13P9YBjdz2uRPhcFiN9inpdGKgoLVvECAMj8H5fdQClr66j1UVlpQ7
5WLLk1kxuhJ+ETqMWhMi6H1pd4wKcJbZVDgmNysgGGDhEiRFtHKzzA4t2XwOclauXu7lkquAC70F
xYRLrWy93ca7tH3X2BNFqQvjNPhgbt4VI9s9HrM047nx5nBwwiiMl8v0qIM0af8hSj0M0jEypgfS
GgOgj/14KVwcmPGldITDVeVoY2G7p5ziRdGNg2RmYb/fnVfT8Jr5Wj3HcOtQzaeGjcvfxRJmfeWj
0NiAoTlzg+ghqpRBDI6l6JFZTN+aLH/h0S5eH35b5/6WUowMDDWvZp+l0LF64sltolnxQdo7WJ6H
XQ2oaLPS3RVGAERS7iEQLABcPgvL2Vxi4vDjrELUnwTXSDHlr7HwlLL0+5HWRJuErnsBs1xlUo31
57Q5uWQtmpXtKVsD0RTD1h3K7qTszb9B3nedF1756ivibDBGgdGnsbHGIiZEaI1EFpxNwIJZrEO2
9uJKp31H6wTuiClQvecxZmjnk1hfu8CEnQdeTqIeadHVFxriT/du8+3lHuIiRSJ1SKlew6cYUltw
/nl82MiL03ZWW8s2ae4PfRkeOg9dXrxSQPU6cSAYwKrR3r+NVyGpGqV4iDEUkDRsmD8l21lTxZKw
54sx3mpDaIgvaSObyFYAVtj4UsU5HTX3S8b47PXxu5Zu15V4foSiZTTGFaKJmvn+CZkRwErJQe3W
FA5IfkLrhaVTUkRc2txwfppjuj4Lr4qbYr4Vlfv5OBfknM8Bu0yfp5w6x52kpBKIKhX3xLjB/ntn
Oi4oCmt5DY2oZp/jXjFi8qERTpu8lJS9buxRygrQdFF2TqoIUyoS2q1GVa+jpBIs8bV5idjIe7kk
/xDEaNlBiygcdK8SZH6YETbyKXYrcqh8YH8qRCfW7GTagWV0jTuBxQmnQTMgU/uW3ettzFt/pDP2
sUcbp14GH/o/VePoKh58esnxuFecpS79tDlCRMmTo1sUKT+bDc9mbiXWOqqXRG21mS6PIOOMus1N
TqqPRdLPFLpozeuOZA2vzmNp4DsCk9LGUJ0rSveMkhLZAMybk/KV61xdhCAWem8Vu07u56sWz7CC
rJXLAKNGlBzMz+lvUTBQP+5DiIYO0X5LBYxy7MH6WC1zv3mk2kJ1DTLDHCa6GzJa+yHElN7ZiHpS
QnPqvdNALDJOnLeMO4iAMt67H3/yeJMys+aljBqVWBwLZ1q16xFiEWFRAPEhJDPQO2XK52ioRDR0
+AhxKzYlTvzEjLOYlK+u08v8sjct/0vxMuqXGi1/SdRsvRFCHvPub0ufPxPCMcKL65A3BNzJx3+H
1sUpKCalUNVsQocDViEUkJxtP9Ei2qf5S9zKZhU+irZOUdgWp6gABPKORUjilXRuS49GEjfXSHws
gpcGU/T3YrlQ0IlFeG5/drs+IbhQeI3eonY3nUXg8xcnOHRX6wK9c9RO1cOyGJ9EgxhjLVJfyOn+
XW+aDTzkaxrwtNtK3RXrmR11JSZ4fE4XGKCNlfSPMTlSf9IZNdnuPt9up7qQRtcgj1LZqih/tpJB
0rQ2fEsD8jvHVRmqJ1pDEbTNLBCF9Wev8CBDg4pU10YR2BTRaORUQ5WO6OoXjXAC7Fe9756J/I4v
WyDq2QceAn769nKX3erQ/uQ9VGTkvnD2u2EQIdDh5zQ8dvzIUFNzhg+a8PMbdro7sRtD5DbNimOD
FHK5W7eVXf5G6DCggew0Gbla0KNMUU3tskiglMAFLZ+RqOc5K78hXQAzy0YzNMquO5engei/Z68j
/8JV6zxQ+1huJEH8OsDDBBdxJegi6DSt2bP9GQWoa2hwr4xf0jX0g+eOg2VxU7fFW8JOabSMa3wR
/1oJWuRwlvycIZYjqpjDcm5xjT/WkqjDYvKiNd68LOIlqqt3GVDTr3AJahOuM29QWuequg/5RaHJ
OPXtYm2D6JBqlKfMOnjdiOCdlqYn1RaDiSTVUPXEzALayKQ0gvrw7qo/GnOrXXAyBXMHGwJ8RXlE
hZOwtfQf8uRYTzEl1J+CvI9t8WXoppEN2nnEFGvzbdksD1VYSCX8LtwaaFUl1tWl2Twdh8KK3Hmm
gnF+374rWWWxgGm1U9OVac4z4/KfIvmOz7M69LbFqCw3e93CcLHR5lZ4xwUasqq4O5ZgdpDd6sHx
yTCfHVc9Aml0St8Wqx4ykqssn5h61id0KxVmhCWKY2FwouiS/8oD3WWg0vrwT84hIaOT57lbuq0C
/rTVvaMaUi6RC8s1GjbBPffz6kGbffF2+WKNRl2iBEEaIJt9koWPu9zDEnH4rlDmQPIsxC8XpTEc
DZY1vZqbietn+NQn+jBNYGmZDN1Mhh/Zuk5o4vDl4BZ6eSBbfLpT6XMVpQA1ugoWRIyI+OZQ5Jar
Uz3/Kbevc5ic+uOFkSRS/LvX+mmQQK6Baud4caiuqrMWMZp8kATRHvPA7xBAQbxWCX3s60SHlh4M
AlKSJmLTKVJ8egWR4p+Biw945FsTqrLkWd+9IFkrf10CsFtGWKSMAxZeIgm3xnRQHcPnqrNzJdKf
9ncnIVHFBcPfFKc7+cCCNj/YRbNIXtP25ctTVA3eVRoEYzQ7EzAU+xDVKp1MXAWUPq4DPFwwYv0S
lBko1Ay1sEH7EghzCx0JTASwokp1Bwp/S79cPZ0FDwIKppSa7fYIImRNtM2nTq2+aJ8nY5slgYk9
dht4K4KQ9YDPWH2PqOwqqYeeNhxmlPMYpbtZiJDVswwTERatjGU6bFcvuXNzNL+V3vYmWg+qbWkS
DG+ZDPTKKA/2KPhKsrqTdNzrpht2eJFI0w21wsY13CciTVzGZXtoW2svEq++9u94nIFT0OO68kTd
RQQFxlGDIL0rsPFnRGFzIxa989wGEnj15v8pYR0dn9QGOXhipBz1+B4SnlkbmpDhs2u2XmGo1USm
qiUc2g0FVvl08pj0P1hkg4S+ray1LJU4w9X3tJzbsEwzqcTeVNCnPAMfMFFjgYvx7gUu/qfOQjel
KjcYKnSc629qF+rGxKTwpU07aZfFsifDASmHtpmrZHgrmk8eCy1RiEht8cuigTQ756b+LEII3i8u
1E0YpFxkUD4txD+OLrmPo2OKQtfUvmuODA8sVUvm/Y9CB9nyjdWm0E27pAN/cisL8jhqCgkBy61P
rGcWUzHnZNzSeD4wB0Q9nZfkA1JZC1nhfr2zojFHqLAZUp2re9WWLPEmISNhUNz2BoCV0IweyNKs
5EE3EDyhVkfPF3gOGkl0d8LN6BbrCGLY4bG8S/bWBPFM6H8wiyxUwLgqcJVz9X0PBoogl0sIJKa4
NXnUYk397piZ7/7I3beq9Ii3A+VSsIgk5yPxsa1FlQll+EYzr2ib6LGVknxBMP4blaJoeXvRW31S
QvJngBHqmXFEZdvuRDP7TRNTubsoELRsme+zc5/VHTd6mblMdxM1eDaoLn5x2LvReOfKg+fSikCQ
E0WcmKqbYRXSywA1A9CEnRuqTwVcvo1vLTNyb1u8ImoqYPYwUJKAhrX4Ysf8LwykgeCmMXHgTdV7
CsRDjMIKwTLp8ART+Gi4Vj+ybmVA/dDLfsxX62OFf4Bj0yLc4QqFEMnXmWVySvNa69XraBCEy4ln
Z/i5WJM6EdnKg+n4AtqPa8HiPIqhNxJlqUAMers0ZXOkzFwlwXj0gPZuBgf9++q6/BWoobqBZvnc
J61NA2/TgRRd3j4McHAjvNILnLfGbk1M3NpsQAWqd7pKd9/NiB9kqOyscHTC2ZDmH7fIvZQzVNLj
kxgk0Lryqg74Tabfn1+XvFVDSlgkYQ67WocLcONwm/QXpqOxRhc5AkpJYutAD2nQvVlZ05zx/Pza
gwBVxjd4VLTwfHAw4JD5pBlit3B5rW3qrO54bZPiFkD+krO5OPCsNb9KmkkewZvR2QV2AACu2cDj
F75gmUgxjH38Mjl0qMP7cC+fxgeHsEGEiurkXyyfmxYTKASFdIKm0edO3sVHXQ5AAm9cYLSF6cNX
YOsyKk9ySooOO9ESSnLmUVC1+cSA7FgNtxemHxzJ7cwo/9BO851BURkI7YlVH7KtKW9MQ9QhvPqF
7PrebWGhYLdcFreB7FO06nJda6eoBPcfABtnfIKaZcCF5d3z2CZN0e3ZoCxR3yzT4RgGYPrXkXA7
O2XgNwI/NhbBiJcX/ZfrbEPKJRlvX4Miea5HykRIZJAml9UqTvQ+1TFKMEaTa2MeRs6YWyf3q3iC
89rordM+J0vDDZONuDXatAJiV7bYJzEMvvKjPysNclMdq5lEvjp8xsYrhcWfUuwLEtcn9wAEUH5t
rvLCPNSMUp0o7t4ID9tNCCL3MEiCJC93A4mH4MmeAcO/8ZuVvXhRraiYNBKHWspzYiTLPiIFiKxr
C6iNA/VLAy3+BY7LGruGEHbItzhsOny2QSMuPfiFFIGCka/RIK1cmKsTKU9kiyxYPlIvflQxlLfU
+PuXM3gDIhC6wMKfr5BZfJOjpmOwWneeC37AfBnLgaXzAHorz88CR+8MCDgwXXAiC+Ck1+qxDAMh
3/DjTGpeNDkh9WgtCYgwLTtyi7LrFaV4kn8N6SepD9SpKt1w89FUiGF4Ijb1Td1JCbV3zIx3GasY
c20MkRDHsd/bQubbaJkb6CwDkRkf3OHPhrDT+iGvGAmngFStMCya8t0LWJDCLkx1a7GwZV0NwCoU
Wl1T6sdWy9J9jenk4O+NdtKofXdcfLOpjTKRediaoQnSj5oaF0Wz3Jok+Zzze2Yup0N9pl8mbLOg
Han9QGX9l87pe+p0ZazjmiFVDMGAJJb86SFt+Nit6ABcXZJw9a3c3AgISz5fLKPgLyNK6TuBp6yE
jEze0QukYlh2e7EFd5E/PIlXtkz7JxqZPWBI8tRARqfOdKyb2c3lSpdJB6F2nMkvet6uRIpVlfMy
OYz9xF1yt0IOWPyYqaMUxCOejxZh6/LCknTNxspmrh86Z1G6q+dP7bPuDjcVEXzulXF6YvpXfSDF
GB2SAx+h6JeF7sVYX/K1imzDRJYF39fkv0U7hy3Au4guHhSH7gZaYZJJgZqjyyWQKBLyGWIkepqM
MVrQI358L6DHz+ZXW335QFn2iq7A4jjrHSwaIStsPjTM6ba1iJNbNZPMdlu1S+BDV8KfE7e0O173
L2hz42H0l203zEB6LwOJIuSjxRurnwjGpr03USs05gf56p9NPCU18gy7hDfQJe9Vw/wMb3wqZsOS
ohFv8593CQQYy7nLHXkwkzxTF/6POQcfxTC4A/FOIvVaPt9DU4W3p2E+3Fa3I90QPM8SrQOGTwhW
YK9mSe4UQ3oEPyIoWoJk0oRrStlvl6MG+DFaKI9KnbkDQWudMdPyEFXRK3bN/JQFE7xO4EB+nQBE
MbVJbTt506NdEr/9eEQWnBfcX3QaeHWRh8qUUPCqs8Hml6SK6hm5U7xANaxrXJ8oOaNyKTIbg6cq
bpl49LouaLX6wh6CkBoPRb/2ddz7mMg6BErSjIr+agz1vNML25P89Zu6l4Q7yhcO+a3nWEJC6osJ
uUKzitBKxuFe2Nr2eLdXryXSwHfkswouj7ONFnZdrS/K6ywWjN9YIi0Z/R/e85v5EBFpK2/iIXTK
a7bCcHX+Wv20xZNjn0n5js9PKS/b4iXab3dkhQ60pM7fKdJ9uZDDgx8psaek8Fc7k4NyEbdg0W3Q
SvVo8D/26LWF6KUyAq1RFWGifxS2ETuRQmLxDTITR3CPmGkHJwpnIajZZ+Z1rTqz8dHT+tujr6US
aRb2lIZTmkTj8+K5FvBvtrmkUUo3X2L3VKsck77jo74EDKEHbhhTBKRd5yhth0vxxdJtqAcc81km
gAY3N0ZXUDakZbuDlQcHMVRvqCB8ooIEl4qMbZKSZEQ2FTS5r+xFkwxZL4AmfNxYLSKiYCD19xqD
VHVKXy2BvCfcCb/gVe/Nvqrm+CJ+PKAWrTd7t0psTOpJm/GcixzrwQ86P3u9xaHJYhm1c7mZTRss
Q+0YB3VIdUo9onkppgTNMVbdVkZxQTGin5OfOR135whNrEUD/zfIfUkz3pxGOk4zMLrQUqBqgG8M
YeL/hCsYnZ58Ez40OWR7EIt6zUDyf4KwXau3UUIy1W5svM3IHc8qLS0N86DhhH5KPHI3JRK6Ur2O
VoRiBLCI9ZL+F36GVBDw4Wq7M30SW3xWGCgp7tY+xEb1e2+vLKOI7FbZKMIH1aAXJqMnHGRkXxSP
SFD5EXaB/eqy0t1ruAaeOGJIA2e1lNldpn04qii0F4xL4SXZHzyjLOeS5lSJn+yRVUxbPvemtWkG
0ZV3JiS01VTXsectlo34B+XOwaFn3ASHar+mzUCijiUSUJLuvFTdtspMlTJ5qBgah2NZzWkUEUNL
2REOoXVmDDkpk7cpwn/fTiK3oBeg7cxUaycibta+3apOcacKjK4yjKZG56TYE5gdQYK0O+qedZLg
D0G7U3DYvMkSI/wGW3lHOVJAwajjeSY8DBFVf9rSQRFaNosLLGQVxeoBllTB88yhr4AKtBIm5RCA
IY1cNlWBnFaYu/+wi1lYkr3/f/QlnqohwNHl57jbEywEbXfQPN7RhB9OV7AuqyH3yscMOgkkD6DI
g9hAG1MltEazLjYO8B5QvDv/5NoJ2Nms6V5kJ3cwzqP9MoNHAD7acq1V9oH0+wICBLNDtr2EJIl7
Pjt0KGX3XfSiKduBeLIpSHuVp/kLZvIrpc+szKNxcPaBCsL2prG2+l5ey3HVEOMLYnbGXIVM1GqX
0Vhqs615s0xgVYWisGpXzeGyLYHFYyQs3dThzjfYcAirbvywlg2Iw3Evt8OQBdRIS34HGa2yUVF0
BEPH88x101RBzaEqjUjzCD48umjC6KMKGGq1DqvnAELlfTrtrNbJ30SHnRviEgC2QP9juekFfskO
/+naYucv/oTHCQbax3TBgsDSJZt9H3iROWK3j01g9PeEwf0YSqSptOWoLBpF7Xl28u6PbCT+NBEE
Z8sLp4uFN9hdqDrPkmOPmmrru2WLWj4iZsbFaLeVbritLLKMAepiIiURcvyNCvbUxLgMVjqzxkZR
ZKImmUjE5Eef3jFCTrG5E53ieKNQpzS83XQ89Vv7vvdM3cKivY3lCGbOAv0FepjzT2R4VQXdVLms
D2hagwiIDJctH+9ZTQMC7MloV/o9BGUXjNJ6U2HlA0X55Hqib+Skc+lKuozbAhPOC4aGNyx+sLU6
aNEB2g9k5gkiBxSOAD1tcj9GFHmPMEsm2zb24FYF74amCBAewo0xE6sC1UG8tBmxWJgzwL8u6bs6
gX+WuWk10YjPII9Rw8o/W/pXtJhmOnWsuBylvgfeupaQIycz47Dw+9XKpvFFT+yd1Xmub0aztVV1
D7KcDzCwyQRrOQUkk2WQGx07l+J7Q4ogJY+tvUFQFXyOx0iHS1vvdGzHYByOA2ws5lRVeoe/Cm6U
Sk5QgVJIpFCW0Pdp9o8xfQJcTf8EamuJQ5n9feo3yHf4ei/roNeFgWvWYpQeKsLMFVSItCZU+wKJ
YmuMfm94zTBj++ZgYU6P6wcS0LKB4vkYnicj5DXvyVYG6jzxifTUOkDqCPyg2CEPkV603Cpimwm7
fsw7CvLEfGkI6m+W8BghqYeCfKLVNqk80fhHiEICVVCffudyi1vbT4K7BX2/H8L6m9zD3C1mP3f+
MKOCrbkmiuIwxCb9WkE3sCGoGkjOG75szWHiXlVrvTYQ4mKOnbwWzOexmfzR7UIYrfVlXj43ZaFo
boCCxK1uCW5D+xxGCLKRpSfKEks5NQj1P/oj9LH+31tzDVWtLfkO8ssmuRUFE3r488oZIbcYy6fV
cgKD+vLf2oVLASm7SR6OsKMb+z5I6TNca1A/1YGstnErMhOq+6W+VB1V/I2KqVXY+/P8o3nA2T37
AWrUEBoSE/uWuE88X65UBNFOuoKnhupVGznUIU/BN1SHEsfdVkrB/h09lDHz9vEowS7gx9iqkjoc
lsYls6RVIExA1FMf4KczurhxYRYCIlVXcn3vIZ7/hHXceyA9Kk38XwJFNJpNtc98nfG3x1sDkcS6
AXKYD514XOg2KMHOr1MSyF31F0W1IoqREgLWHurlIF8qpEgTmL7pK3PmKF5ILr/zEiu8FGAg8V1l
WV29niQTnC5dEuT+zFMgjSNpZj+dmeoYXVzoB8rGOaYknWWIMtgjefjwXJrEScqvE9Ru38Pnkm/u
RJEy9dPc+CiTG29IfahLqr1soSazuK5uFhd/5guFr+bKmb8FMBTPVPESjqcv4rG4oa4Se9rP6wfW
evIp/FpV0vqLwYr9l7XkLs3iPo9owErNeyuSovYyvAav66EmlPPZclXVd2Ps0Udnm/an+KJLQgIp
yRWltFVUgRnQoutwzBKDG67xnfzzOFPcIl8ZFGmLVQ7L3pBLHaDiScshWUMqjLENP5spAZCfUrjo
opNGwVPFBkVCUU3i0XPnlt8V9j6zjMT20sUeQ7k9TIByHw8rYhuxR+spAF4iwmwuIxXTH6BgQhF1
QyINdjtezScERdJ090MuVTYSDfMMxdCLduGxukrp0fyFxbftJI27GiozdE4CsW9fQPhNB8YQR+su
12jOmHL/ASA5nbj3FtmxPLwOYF90CHPxSpZD4BGiRYIyf37RXkMZDekopzeHfoPYqdPbyjHLwl+H
Qg2gZy+D1H4dmzZRAScZclyC0FIqIqrKm+hUaycOKbCWR5m5LUBQEH1AR5sMfSlzBBaR+wPIHPsw
wGoyeuF1J8i18DDV6XEVLQPwE6d6Df+8DC0f4KtO/3dMNvxwIkZfA1mu722sTadbcog/61xYotWD
xx1oI4Qa4D2CcdVGxSgI6vqYyC86c6TYIuNbnYQlJnr00FHaNyT/LxxxkcU2ni0IWR+Ix4MiVqIL
VYH7h9DtCePBkcnFq7FykBMZ+5o67cnedFUBL7ywyx9waJ7tSmjXDyCFQx6CpL3e30v5b5BP//RX
IIuJsKT01aRnbe22lLlxPLbAuRXB+BW0QQEwMo1zPVkv/x87HkrEIx/O9ncjkqyQNuuXASWeJdGS
1J8N/382uyyj+1j03aN9mGBGf5b51UcoHC4yTkePzHa/p106OG+FgL6bF0RPBWDkwnASjIxl0wLt
Kz7Sf8ZkTKrDYP02trKn1mBOb+MqHG+ErZpNHIXRXb+0GFjZay27Jx2iamXgtKWJYFkxux3l67Yy
YF+9AxFrVsG8ksnJa6LhorBj6q8kC5vqdQMbEYkn/+poXaMfh9/ZpHHkxsddEGYyodeoF/7odHpZ
eUAC+KOI5jctoUYwA/uE5Amg9XfKkNLmq0BvLOk/vdf8FF2TtATBUwiGGBNbMmy1uXDOPeyc9aHn
bJK6VOs334ArH5OP12ucqDoWMalC5I81SwpPJUpg37xh1QpwJbigpyt3TyElZNeKx5MVyljT4kL+
YCh/onxhp1U/o84J1m+Yi5ChdL4Fx/JvU7mh6olx5luRH5k8pk+64N4I6CS2SZIrUlLmNTqYd+I5
WwoCPzJDuhU6rfFkFwk6cbeqBFnWQ24y72CO3EGRVIiza10WF8Pa/hj9RnAmLMlVmQD24mpSGWYF
c9ZjwftMlztXW86J3kSqvqeQ9byvBtBkh24fEM3SrmRPGYa/9rwvNGzHC1BxPBwUczyiyCTEFvIo
sMmeEae8v9xeo9gtMFJy+gYx3HcpwWDcayGIRSp3FS6SNRCyh+ZD++9QMNhaVB9K+yDd3HP2ZunK
ENfwb0u/arFq8jfzuK+EzY8//fmExZTWFphDkzqZg1am2qFOW9yZyEbzxXrwCn0el1bzST3vlsy7
PDG9xTrfjECUP4cw1c3ZmS79ehNxIbmdlksV3t7+kyzebuuB+aP8sr3MR5kUOP0NPnXQWiz/Vop/
sbO4EoeXvcy0cwbWcJlU6utSSC/5zqhhjy9sx5HnrEt6cqG3128DDgPEVQsdnAB8mGVeAOUghqJD
UaJIjA36dQHqFemcVqzAR6zolIQkNsdHU32EW+13HdA2m/BORbTsgJJ7Evtm2vS5Oml4+4T4PsEZ
Nmnz0X2VcTG8V/oc6TgksXJoeWhytKBwDGqt2eZV0CvGmg9oxCFxDLYDSdlOjeKQeGVr5AX+NqZY
Pt2yof0VOlZlYWwW68gvtNhh1nkteYfh31RoyOvxWx3fsrvJZfcl1lO+a2DoJSY6T/Yccva3VZbv
byX/2hH5BYH2r4dAOeCgBiA7yo5QlK8fZmNzLZOjKJYhVIMeXU2xIFNeCUewDdlMhHFv3WlNV5hd
gFEB7azakrUnGMuzSMPgpFmiKWGD/rxV7FHpOzQze3G6HNxuAKlihw92ScbgUseJsB0K42PUdwgO
bw8ck8yC/XNo2wTuwl76kQpYfg/yj87nDT/nZw0Sy52OBUWoypZyBejMS6LVScKr4rEn1XXA99rF
B0FjKyREUHGHzK117wZkAIMfu2534bigpMiAHo6F7wYug2u4uZDx94hUMODolFvQCTlOkFNXz+zI
dMNrgCaSC8CCMFvx9VIQQvWHRosL5r+qJL6nKLBgpE4n9mlfan9j87hixEllWMutazYIvp+YyymB
FeKuf6qDYDDIpP5EkccowhV7ZN6+xFepslMXRvYWv/6lfx6QGMzjumuf+AmigL46Ly0JRILSiXh0
4UjZ9UXLeAkV967jrRrWtNi+w9NBFwV35Q4G3oxEEsEbdc0qXGXZbDe5kiKIdi8pQUhzjMIbdcgw
eGn9cxnZh0s/BnuHX92I6FWYqaC39RB7jeJcyNzmi6m/09UVA43TtBJQuSitK0UGjS9sRpxYE8Fv
iYPMDI3h5/ulNpUwL4UKf+kIF/QbQuSr/ia5u4INPEuztzFZ6KN1EAvlZcvH5C3K7qWYmYyXvDbm
hjPD5MVgAWeLPMihADV/Y+n3pXU19lZEflGwutJyorPYrNiDZJFd/SmhIZAc0TZA06Yp478ydLge
wGPnFWUjt9IhtZNt6GeuWGK/tpUCBj1j0RuZXkUlem4BuLLgGCiM9JyhsOAeDB8aluSfX3f3W3qZ
dQxKCKgcj1JJrNwFofn22e8ZfQgxxU4zlhrhSk+ji9N8WJAbi5fW/hg+7WlRuBf4C5U5tn63TiFX
J0xJC+cT3nJkNYDVLxhNXPqOuQfr19bqVIe9ByYsBR4E0ToKSUIp50ANma5GAvytyK3ayDGNnMYB
RndB/q6EreASarHw9Mv3QrOCND2MLQOvAGp7QFMyzoe8OHoR2FgEY/XY3J5pEzomWoJ+jGcPVSCe
Y1Ns47V0fSOm4LCf9r13ZFm901d85UWRK/xijP5BwEMwxLHp9U3zQGJTQj4CbcKqVubZY2uka11V
bbteIQuEpGrV8SbJNxDiNCa4nIig5rUmEFpAfyxGxelz5FfFv9LbvaCwXsM0zAjCCFaury1qhf49
6B4xH+SAQP4BVI9o5hRJrphNxINqFP9+h+s1keDQFCfRQkPxNShTOb41JFR9BverDT8zrsXz0Fny
oKDqcf909BQZFnhbA4xo8KINP4W4hj8J7Y0DCw9cLKuhapzw2DLQ4Jx/38wfGtH0BpbM2ktO/AUn
IDuq0RYnu18GZ6Z48EEBkKvNJKj79MyL+jRqjd2FoIaT7RQ3uBT9G0h1+DI97bT3kFIVCtudksNA
CfS3aPT37b/1dgzrYByMZy3TRbVwMtvqjF29gsJ7rh2nHjZ8svis8qztP9tiYo46prCwfVFCNbJB
YUoZmF9K4J+b0yXBA9uKV7qTWBGEekgoGFThnDbljjt5vCqSsv0sHu/Cvi8qYb6pwht3Tj+YzWyc
/lg18MQI64BOAyvUpzL7/7Yi/QJTGrflstAx5H13enOSDzbwJS8rPh8xqb71/JDqDDu75PESlNzb
rBZy5NCGN9UkJVPu2NKGYZF2PAzSSa0AU1lvdQBKZFjijRv3n+gqXG2kEAdlRPULwVfvfc1peQPP
foEApkuACvf6r4LSSt5FmYYHctNNhQX+SzfLOviKJN9wjpAE5qiY3StXD/q9X007478C036r0eUh
sGb+pNzBfslTlv0USZlyVuvoENs64x1X8ZDC4GU+vfmEX9O+lSY2aWsr69IGlqmFTx0TIz1rzoJq
lBwub9bVOYqUV8PXT5cvpY0ojycApp9FCJk+9ajf8QMKrIw4+Q4pxbClTl7M1JgfvnRHk2x2JJ3j
FKeaWaYw0+u2ZPrM48PIYgVTcWnhKJ0sPRUYuAj5b0qCqbYd3LCJaJkz9mpXcv0WTC5PyUQr02mc
bJjiXQBkkM1foRM9G/3d470QjA+ZihW5ntv52tiGICjOqftPA74GRJpYuchnOHV0ZapqA222LrpO
Hw+YZop8AuuXfwEEgmpf8qJptFDT6xFrtUGFIVY78JP7aErKoBI5lmTFLH8d9ZcEL7lYDtdIHLhM
5TSrceDn405d/qt8Ojth97zYvEgHh4uZrMHaThAqM216jwGR8ZA1BsbHY0bLw+9HplLMIr8UmNiW
VULXFSoecLmQTEDpkrJuGVhegsozw1SiHt+Si3wUAoxVbwQKjqLvvbi6nHm01Nr2Ws81av1UUCYM
isYlpO/gsz5z9Rj4Rw9aTQTin3ucEpmQfgb5VB+sDFU8HGwgnSl3GjzTqYXeos6EpLJ1yOwtsvfb
v484EU24uc4G28+QNdrIEKAatXR7NU6bvdIjt66jhoNaMOsxk2z56HckLIieAe4TSPOd1eb04/GC
/1gGY112SYuhV2q7cHCdco+2UmR2KO2G6GRFxUNuXW72VWnnrSX9ARCtgWsL/mloSv4qwBo/Qhcx
oh2VA8Eu3HGZ5HuyqxX7QEvbReHD/xYsX6cxOnkR2Qz9QbYW+D9xxi+VgPam3aUCCpfhR2oBW/KH
YOtZeLiieEAlG8apLdPVzdY0B5+RUj3iKp+AMHCMtXZ/5EGh+51QBSlWB6SzuVzgkCY8u2aPVn5I
CVYoevcQZuv+edfwb/rv7/z4iUSeHbv3iu2FUKFZAkftRMwcwIyH5XcBTSVFnTmcT4Wzh2W+7i7i
yKLBUE1T6Hd+kb4BvcQrrWvhkWjG6uNgvhMdO8tCe/QVQORxefKXEXsatfQ5wHTIaqR2EiuDEuUe
P7uYMvcSuKLFwqp04TtIRpbjaCpJJy/Bo9CSgPyT/D12lCVhwj6dO3d+rUJVXPFFeqkT/V/69ywd
eALjbCrBezOm2y6DbbE2HRMICsZWtCxPDVngm9Q4u/FjSWVvXccWySe8F6cyK6lCxSVGSwmjECTh
V7PKbLMwxAuddI8OujTqvEFvH3FZHv8NRG4S3D0n3uvfZjjwgJjF+dmEzNFivpjF1saRZfTBHmG6
nuIZ/fnKhwzvZPkbQAfwdfOBZZC1GB91O4tnc3IBADbt4f/Du4YM2xV6X+W7y836u860p/p1A8Y5
+XR9isvLxOouqFI3gaVFboWL05NTAx3u08yR1NOirJXIBfGQrzT9S8BzMYhKYc4mbs1Pyaket2X1
TCOMWbHRkmWyn/O8sqXRxZM+aD2GcpH6s5DmWou5NBqCS9oy+s20578fKVQ5B6+rawuxJXdvXCpK
vFLX5IXmipVhI6id+MjM+71ce5LNwcDMTX08mcbV1+oe1EFYctYEiPg8Z48C7oNXeizOq0VTonZl
R3J6bF0GUpBikc2qFRNZL9XgtgfThMjzb/G8td1ieCx+bYnD+lRRuhT9vIksO4yjnqBf77J4XULr
AIEvxMnfMyVURMrX0NxTRZDNFN93M6TPzR6K3xWC/1x4trKkLHXJxE2ZuaA/pHxcSUvVyeso7LbN
ddv0p5WSeViG2adD2C6lJ4YuKbXOfT8LuhW1G73ITdvab0e+yrmaVb2AjHoI3yj9zVfBJUldtbnk
qhdyPJ6iT8dX94benRl9Vakfc3wmZQRiMHiVjPAGGtY8uW1BBAjjswQHFRl3I3SEjAEBY3oWeghw
+NTxsLEeGi3v9rmOIeENZwWV8Ht2YgYiRto2FBEMfUgcHznFWKJsGkZAiGpuaz2j2RCzxfgJZdkN
WFAT4Atlry08rJtYCNEwjnHaLW9R3HPh1aVV+T+h6QVX2Wie6RET3yEa7XxWQdlBQLa1iBOx3YoT
nJCnxSPDW+qAwFIgDx50GFi9d3NyZxh/Whw6FpCHuEOXlx6ONB1AtTnBetiPwIbgcXECIySd14nf
j7canCOv8qg+C0Oe9b8jrGPDUnm1+eipi6Z4S89HvNbuKJ5cAOVHCM0xGeEiQRfWdDlNuKHoelnl
GbKAFAB/5ZwNMuQe9mey4JOMdPoWNbEOvHlr6yyubEtniuvYPseJsShf31+aeBO3KKsQKUzoqq45
soJHANlntXc5/cd/wx+i1FMXwQwsU5MNGJJrvForPIMyrYMXpRhuN9HG6SaKaYSG5luwFF27/1nS
WzL7Ygbl82YLdu/Uv7FDnqC3MI3JvNjIuCUxBuwYnUDSzbFi4Teoaf7yNddSJbFVKSFK4/23juyY
MpxyXSLH5esHfEu1IiJ949QmFdhatSh0x8/BCvzmKOQHcPu8EXpfOrO/3pdwYBilSJ88KUrSQqIU
pQCudLleFwfAYO0mDmj/cXl5MeYNW8bGBGFDtdEYHRRq0MQlM+DcjaRtNtkhQCVzaaUPhCf7CJC0
k7Em4SIQL+boicDZu6Q+EseCClzHbtyKKvRHwALrKlo1yz+6/T2AbBYxSeuxdRGQSdtY17WMljd5
8gLA3b5W+D+nywjHK4HkbFxfHOXElBZohijqD7t6FsGk1DNXkBQPBfRKld/RqnHMONCmACC7GKiL
7fPPVqd7Gmh2Rk+Aat1FZooe55bKwuSwQiM49eeMK9pxwDdAaAxCAbp2AOUggEXbOsM0a2ItUORT
koaChMEPsIoM9xWn1nJh2mnrKgNA/HGCx+vndw5teoG2gTeFzNd8V+MT5wNd9xCYoDsIxQzOQZNm
8PQOOkXZDkVpwPwzJYtgYdHBLroXiY7+4d2UcQ1KgtfvVIbned7QOqsmq0LyIicU2iH7EHy0/mAw
0fuS8hmi/1gEF5JikK33GTGyx3j5XA5ztfhGKP/ZFj0RipIsM7D6ivqqVr4tPw4DbkmwYt+M5Uwz
21a9ecSOYRpNdRFPuN8xF/Xbi21pyn9NB48hO5a4NLUbfKD+hkF7GIx0LK0biXNS576kA8evJlxg
VWtAA/ZbgeurGEAheCruddZFgri/7JdtZrm7RrKEThZz6H/S4JD61g86ZMqHsbLHnJtSEtc/YnzO
C6mdOROtd+0HVnUFuFN8BnwxMlJA6jmOLPD77uHc4T0TtZrzoy4oy7HK3HfdGXySfkDIQQL4tjXA
Ynebt81DW96FrSD/S7hMyW4mQr0dAGH0/4J3TyqYLhbpYN4cvBMNuSjK9+w7J7PTbDLEUMx8/k3f
K+ZLg0sGLni08B1eYy2inEPWyuX0z0K0SJ0Q7bGU7RpTXGdf5Mw/d1T1l/jKQZyPWTID4sf0J2m4
8Yz69/8bdsuSyJ0ICkGA01l1+HaUTNMj0VQpkV6zZFzYo5cP4kTVfpXCI2rzA8mlMVTtn6MYRJND
fPyU6fLQ/PXT7Nnrt8v9QV3f3VDRZpBI9Ut9rKGoRDra7+la+ZcA+x1rM4jkxO2kJSuBXph2ccxp
1pBGB9133QAhu7VuagcR9Ef/Ng/iXn3Gc2qK7K653p/9G0ERKBdXeum7Gv1jL+tjIDXbihK8JgsM
4IyTil3odtLjMkgP64goInnRSiMH+8Amyk5Bm0uh6v/buNbne12mgUsvjtrGuRmW+PBUFD0Nw9jj
ZCUlzJw2ZgilRi5s5LgaO2t/us44uUrfim75DSNL5R8RtVrA5K29snaezG4zOTWnPM+MnzRrbeT+
V+z4uz4hjMAC2uc08S8M5BXzukPH4ago9iPav3vBHvg4IG67+vw0GETM1Xa7sldvShOrBFUeqqbK
XDCqLyuK7bkjX74vtWlC0lsNJLQdONr7bDOsfadhS0EUoVUL03QmZJl23kKYMVNvy3/dQlnXYT9I
B/XGhGVhQZOe358fVkHon1JplfViPmpiMdtN1yKwwEIYX2qng+KkPInc79QJ5MAzMrbYlhoE2Kkj
ZcUDczfKPTQLSuATvCstRZsmDo6HvMafxtP5gdLgh2lUoKcsm4agdnF/8kR+iCxr4MhdXw1LRklE
vmc7AdT++SjjpeUvFOqwSQtttcOIrJq0Jn1cjGk23VI8KzyeJUASFrAXLvetqmthFPbUIAV2zS9U
hOAYMAS3uNFK8FdvJSfPQLrJ2P6gyETN/6HmDSFXO9gVw4ktBJuOu1sMgMsIQ4dMxyjDHm4HoRZW
I79SDgAj9Rcwp08CxSd+kvGcCMx/7ezwYF47vJzJgPzp774wugln7oc7+zgYZl83Jsw+2RoDE/wn
Ur9mNjpfjyfTiCjnLf2+8xSnLzsbEwl8N9PmuY9ipiqSxr3HAr2MuieKZVbvWgnLcsMaraXiuwPL
w+PskZz3vZgXJk/1QkTvKM3xVGYgbAZtztZTAVYcyDL6jTkyFHksZA/CoxYXH4i+DVgl7NelMZCQ
wt9WRlR6mea6b3pnqozp3UKn76ByL8hsBUu6eISQPO4jFn7/+Yo81IOhCK6vpYVPtyrZ0v65pdZC
l4+EdpbGksgvYzYZAp7JEh8jV4CJG8FrcrXjnE45KRIcwn6V1OyRfj9leIJ/bF8KzpBfXc1E+g5e
qiJiwdWXkkcjcDxqw2IfaFlUBp2o3uTOsRW9FU/4OKj6C6gFoGo+cFxF/XGCa1V1SRQpGE/Pkinr
HkSMR6DDbfLmZOThNQRZapnYDWFc8A6stbMtI+eJVLmKC9Jlg/cZGSiTpMeMX+DdJLEQAOU84EEM
hyTxwVsO4mdYw1Nrd7hctHpviTfRgO+WzBzCDoBZ4KZG9ToYvUtg+/owPWP2uGNXnK3bvevElHYw
Karw1X9YtwybnLwM3xFB+Ya7xFZAJqYdyMUJMiEDiaOWIqGc1XX/TYVPNtgUGCRcvPx8J7ENC1N3
/aJrqwfhTb+nhlLKhx4VZhGuHvi6QIsQC68M37RA5UyNYRnhHDMir1ryI1/Ahml2Lwua7nu5STOr
mkm+LcNzBweRdmLsj+j8vPVvqr9X0BE5msQz8u31C5pAe58DvuwqdWQsASQ0a8YJVrgNmMzszffG
Y1y/Ys2g5320ojEfsAlqfSdDUaZ/uOBEoyz39X7kTUlFN4QsLI6i+xfR930rT/F3plMj0qI9+NSX
JJcaDirMMnt40l9hFKqAhh+k3O/DFuIOxGMPppzNQWsmSeoD7Gm5bRokGEzurMULyRJCVTXkSsUG
Ooe1l3D5iYRybykuXdtDLLEaTBKk2IAInfJuhNL0TLOeyRarfrrKJnXUYRv3GbOYchmZ1dnbVXku
hvWN6ChDqlXiB+O8E2fxsxoGlbBMVK7rspKK0ItJpFrlCuvmNRLBZ4bmWyxMMVcpPy80uJYM5oF1
iAP7BAIKdnNUesxrRM77JcPIk6nHOEoLrJQbJK7a2MyZ/S5D0qqj7OMaVja30U/NDlpIiys9l4sS
oqN6LO6wxK+NLqTN0FHzyTyH97CKQsiqZZEvIJSz7/bzcYJ8O8G4vRPdLfaR1Bn+/7WlDSgkx0JC
U8hfFIO4mPADu4m6ca4D8NhZV3+9mcgamr6iDkl3CkY/1jg4vmUrhR0DYO2bB0ZRyPb/mWUwvuyj
PQbSsYhCxFhMR4sEBKxCdefc+N9NeSHN0NbA7crR3cfLOS7Lza/BzH1ypiDtn0spD7HoHb6ACbYM
Gejyh2PNtQgI2SemSyErObYabYtQIeOVCWp3hr7QeC6hDmVvPXcfkxUpanrk/UektWVYzEeCcj7v
v5w2nPXHQ12ulcoS1PTEgeds5iQHQDUdqX/bXi2pkcdptnLCFohz3o/haqmOUWGbBVHNFu9t6Qs6
3qeXD+chldPP8E0MLAHfLFcRevPslq7oKsZo1VMNPvgs3m+jOxxhX5oKtsmxfMBdzdDhW9w0gmdg
fDgBFhKGuom7y+vSN0k5uZAirn5mgK3UOHw+2E+5gmFN9DARNOUXCwZy1bb5E91aQufhhLr6OQhi
Ux6XvlCTCPY/CoOFbdVZ8ohj9SOZcdztBk2m2ndBO2/5X+oHdDyr0ifCRdItXZk3tyiUH93YxzvS
bazK9I5G5XKS6Xcy1p3yPe7jgZK36mSDTnuRg/ke764ho13GeULeWqJ5rAdbTUmzKblaF3eNEvsk
c8YZvEd9IdZdlgiIQ9Z1epkDNoXx6c4iErbK+DFS8EEVna3Lvo0PhrzArg/+qOv4FuHP+Nbivmvb
/v02aOrC/M81wzz/vaZCfa8dwOZDv0pn4FfekXo36foHA4RUQRRaAHl1+wTnUvNYUaaZMNMgn9/D
ocOlt8sElxrT7ezln5n2ijQ6amVbZy20mqCmfOY+CbwawOV7NMC9tyG9BzidvoramQ+Rku30uwK6
XPE4kkge1EYYkxSnOG2iRoj+7DJ0RQpk9ZqsLZcixx8OFsvvmTRv2pOh3MZXkE/niH/UVqHNjebj
taKcx+wRl9EiVnV/m/Qq2u1sZLXNaQnS+cMXn9TRjCm+SFQQ/n32SM2o5ahdlOEqq3YhDNKd4Emf
02TNGgu+KuPrMckbdtHn9/+S1nhP9MLgx+vNvtoMkKNRYFb/gdQzMl0+4QyHl2rFTaOLbM6UWfFj
pepvwp9Qjko+DsaE3A5t3SbiUta7Fyg62651KX45zydfQ7aYUK/YQjn5zRF6K3idkY6sPEHCWQBV
gN7ewvXeGBHAlwkkY28Fqjp15xq2puJsr58lhf0iCOXyju2MjVME6g9TLxwucrQ1Rhz3/qmxp1YA
8B84R9bytAyH/1bsq8u4s+6Ur5Ih1OvW6T8+uFpLVHL5JSZTCViADgmTKkHON1Vr0/lnPbWHsed6
JZNUda+V68niWSE5e/cUUF4W7pu/OV6Lz55qxwY7kU7OC1d2j803mX8JCohevHeLOhh27dz712b4
t/UjlA3HyJ5VYCUThlQBDhnptJNxkqBvpppXw+kfzGESqh3T7FLXXfWxfenzLzXlNIEA5oRtyb6X
CsHS0ACGifNdDI01NhA6AgewArSSZVWtkfwF9zFNXyZRkUXl1aoO/i78dGv1Jvt1oR/OVhxnvDCP
c6CYLQnLC2jgJr8EwFIWkD9j8O20ZYUBUs9MXI+8anFOsbgi2Mu5BYvhpunOMbaR6MVoOpnFjj0Z
neGdQ5HVmYljmZfgtpF3Aqs6CksUG510Qr8jv8H2rK5ah+BevbrS/f6y45EIG51HfsAMRNmg4S2g
OJOZupipnT00rwev548DzRNPSGyrr/+hv8p2mv2rdOpjlV98lRQVxDVVD9TGQAXZKh223oMy9ud1
jllLq18rZ/JppRfV67Fyye3NV7bnZyGygvLzbuePu5r1fjh1SlfhwGUvdDdw235xFuf4Q2o/DTcb
y74MZziRT2aEnRkuvWQTaqBrgWDyejflIBvv+e4zl5nNC+VPGjII2Vqmrb8nSu3OU+I1JhWYg6Cr
MFOpLQcFzOBz7uX+oaFlwjtOrBrBGyl3ORf6PAFPYEA2nh8u1Ymd8MW5I05urVjCoG6xZPLB+whW
fnOoSGYd9Vco5G+sx4Zaf2YBNr4z8wKs9k4qsvYNk5ZqITu3xdFlITe/JtvqQwbDCrH94iwocryu
lUzSfMfCG/GBTh0TTbOFQWy8hZsBxhP19usXx0vjMNCq4hUS/FhUSd/n9m6P0nzDVCyBmSwufAXD
0vYTOgDLSMn8ymyvyLVoUKN6vmb3wZKArzklJ5bg/um0c8qXrkqArEEqQ5RKDg0oq7EhxsA+yoWK
tR2QLR62DTiQ+TkMvqUAVOhT0YsU4hcx0X7U4w67eSB7+1Gq73aIXXAeYs7kL4leafi8M/pf34WD
csggguHYGOQXwkZ0B2iGOYga7gmuzHcrVPSI4ZaENRpDX4AvypYQtKIGjXT+EV+OYZzK8HDp9w0R
IFecGDKvuLEYx9PzbC8HiWZ49jfRSZ63y5LXb4jjeb5tqcB9a8Zc447NeWGJ/JVIcaazu6ECqvmN
hxn6wzOYITzelWSlfIFJPhboBoqUCC52/vQJm3iXpVtoTzBwenqaKp6xC5vlorZfbH7yPe1QhY7S
3cIJlqEVenfNwGe8vtynHLdqjEhEdbn5NVzckJxkdkZVfleLVusndTomuibB1d64WZjSBUu34AOc
Tcx2NaEsY24KDAYvZp8DuyRuNe/kNyLqGtGkevuBZpG9vcKr/xUVhYK6fo5N2ySGMe3Nizy0qmth
xYnwS5/Jbm4Lftql2Y31Jck43hjcqzhRAxP0U6HMvrUi9UvpMulo3iSJPzVehME+O1mUqnYgwXi1
ZqF4BrDYW/EVLvwj+jEwMRaklFASDj7wQT1zsvmAETKnKTNXXFp0QJjrXbe2x+q4emtOf/Rouda8
X1Dh93HiOThHxNgorfdjEQqTWhzh0Ys+Xp+Itkmnw0izx47C/Ow8VrB0OzQ2KwDqVxMb8jRaS3zp
zXXlhffbqXDGjYOMC04+C05zKiUu+uGwuZd6k5/HmgQBGbdy91fZgTveYK+KVxh0B3uZaBfdlkQN
1FvrorwJuBfOBq9+jyjzCfW9jazN1Q2f97UM4GbgED1yhbwmmy9VlcBAQmgjZ0MgqwYE6yUjfCL0
BeHQZkSAtGtQp+jjdRayMnAg4JWe4u9qxaKSADaMFNwmtgIsjSGgtd6XHtULxC5XIdO08T6I8D4I
6fL6H09fOQWWMxPSNaq52Yw9QcBZAPmBN3q1NVvXnajkpFjOE7djRLCPxbaUQFMqNh/qEuPuHjP7
mADBBTDUa7hcylV4uC9ZnnsMT5UnzAPOStsbcRLFBjyu4LWwXCJdBVtwyGJgwrv7tpA3R07wiaMa
bfuHQH9aqcAj+PEvfxi7Xs2g02jevXfu7f2jkscCt/i+lZutnMxM3EwNIzD0Tt181dHmyoiRe4b4
6p0l5bUqroeHNtcHIOotEiO/eW29N2/wpI6SvgBGeuD5fkrCPFkmseXXUVv+JWe1MH9OajgFQfb1
opzmF3iy4LYd+1yeNb/sWwC1B4iYHryUvv6veoiRnYL0Y/MaChP6XnyXi3KUJQkLzVtkGNJa1ZPt
0zPUd3SVNEYSEgxTip7iqeiv1s5LgcljcXPpZ9OsQbEgq01oOaoPCQYfurivjSpl0aAMHZUpGJjk
YO1ZZ6temCHyzfEAOuSC8S9SX3PyOEfQGb34NEZx+y9PsHlM7QdjOaSUhl9CpOG8MV8Ld2RXET3t
7GxFBxsYXJFjVv2xtz5Uz2kfjNN7dbeCGSCWG/dbLX/38ZWbhNK5cO8ZNTEpGdZuMeIEWdtUM7PH
88C37bwvKB3hTzs7AHsremhlbJC7W/oX5gooPwKms1D09Tqx36J64vh2ZmfxRlGd6lvOsgEDY5La
77WC8iZPg1g/zViBpAYmr5MFjcPim8Rww5oQtGdM9WmSteuIaEyRmapsTADOFiAG5z4DYwOQbvbs
ISBfiwJNzZKKfMrVAkCtIq8hiI3aGVONFL+EZUh2qqHSlVVwU515wc1VjNGxZWJb7o50TWls9iSy
BsNrqmimc0E9MgxCNgplDVe1DkeF6bPVlE5A8to8PkIOI7EHERMPQSKFdAXtTBK44AQ00C+wrRW2
rmVN8hPyddgv6yhWRKzoQBvD9/Cf5KkP9ea+IsTiX/EV8thIsy6qRp2qFJtK4fBEnrIU7DzuJEJM
0/Zf+b7Il0hrJ+GKKqWvfi0z6K+wy00bXIjwXdSAxuriceRyXGh6LlibSCqZZLgKVoh2EMNtr0AN
qLx4sYl0fJM8d8QI7lbTXy4qEdA36k4Hq59BKybozZ+edkLogku+9qh5jTN3oEYbYtfTWgwNrpHD
CwYbwn0awsFzp+LluRY9wvCMa3+PW24v+FBO90U8fvHHCN/+JY8Jzs8oOt1Do4AT7MvtIqel0ovE
PrW+f8cd6zGWpoRh+zvxGXTF61EyPHAxVK2pzSWmO22xMHErltCLqhEgxGKfMp9oHTIZJS8akjzB
2XH+h9sS4NRhhLPzqc0PhisKib+rkvk6ix7jmI7CRC/SffZJDFKfn/NzMISzNrk7ES27ZaHViIs5
Lv1Ws0UUn+nMH2pRfx6pp2ZVtud6rPVUceIvJ2wwYzWPbBOT+Z0/t+1ha2aW6QtF2hCV+o40qMsS
B5nNp8bcZU9CXWnRF0MQd6N6JK3ieYnG4/SPpMaUcI/ZShHGFU+dN/sI7E04yI1x4BzjULIHtYzC
2ciI9yzwEfKJ1YDlree2+Jv7ErPVT7cvAfHe303gM70MLFPy49Kkcq3NsFifAuU9Ys8EoapljZL/
YG/5fa8nzPZ0vicJM14RLcEJoRbDA3t6ULxtoAT6ChWoA5fHUkczNndOdNcqaLLsodDNZfqm1D8v
6Oxefrlc0RF+723beCu24ZTwadJV2czWOKCqKaPHVCDGKBA8SddYB+af/sWwaqzkjY+zWDGH1tlx
b1aOj9gqpEofkrlwcrv+6rN9vc9VkBVm5/NXyxo2O46gbGrYKybL3VCTmFoimHHIkGaNvf9T8fko
1Kz7GsDrz+ldSpZltXq0B/PZUeVGyUuGGZbNIS3qCLTymGX+yvZrtbo4qlHg7/9asCBn6VWjePjz
4/eXm3YADQya7XAzQn6uXtxcbJCSBY6BaknechtUAtaa0/bIXZwJw0ske1NsHS4zxNRmXVJvDj3K
FdGhTqlL90N/1ZMeNekhGR2s07T8vcxEBxmS5TiIGkK5OwjVNmjDiuvwx8oDJVbVmmdIC4rcRVUl
x3kh7exz3e5Kaa3B177wbs/MOuFj183XM+TH50jnWn6aqaQMqAs5u5aJqH0RGVz4n++shjZ2Mm/r
NodEmQ8mHX/z0aD2wXKhJTRg9wGvy8cst6Dc4nlYzDLBY47bymaddASFzMTUsWXfly3RqIDg1jfn
qIaBll+SsL03P4kuW+wwxHufQikUpvI2S/FkYtdOidF0owzFnlsQY5VauQ8ss99yyHeMV3W24C0d
B2Pq0dbrjGdlU4nIvaIS8KdC/wO8M3QN88k9mUTMShBTXmjA8xp6HXAWC3bTiE4pet8q06FqXEDI
ZaqxeBYxssj+g7HI3nMvt9GUpFNb0PFXa7TdKq5JV1z6FQu1XEMvT5Jva9PD0YeyV/3h9eZ9aa9D
MhgM3KevMmYNUCIHe+S3P5m8ZjJlxmQTLo0FAVKFIJ0C/fusnJM0ahm3wAJJMk0LLaucOr0AMzC/
dEU7l2MygfQcR+YpAiKScCAZW6YzIfjHz2RcXEvXYjcqBg2UrvQfzE7dUm8lPf6NA1yrQN9LGdUM
9jmmZC4xHzXvzghRx5hKupK5LyeQfS6Ivpze5K/tSK0ha9n/2iQPaB4NJslGjPpqx57mo0zmsoqF
WgrZmsX09G2gLOCmjh0PgQtKragttkUoyz30ts8nu75ua4N30xiJzKgzyRAO/wqWQRrHZ49CUGKy
9P4i9l/UZ/0Q8hv9eU6cZsNL934BlhTxMh67rT40vnFBbbaeFJKDVPlMUTx50jZiDxyg9qy0ZMLY
2mnRhwUTxEHiKpYVK5PM0aszNxxkeZC+aVk9PzooHRbcJRUOtNuOgEjOWuTAyOluF2k8aHejXtjG
zZL3VGMHIRqG4XFqUiuASBBznRZPpS9fzgkKj2WjbL6SNTgR3xB1J6Zq20j1NZTe41/Rt6HeLapM
aNq5NYJXpS4XYA+b3Gromo+P2JWM0njaoJeEyb9Pu98eknT/EzrXipz062hnITFhy+l+SHRsD6t4
XQRXgdVkPdJTiciflGzijFLq/Lru1ZeGnvOtToT4WXOAmeqH0txJ9ilHpUIpC+dYU7/ELJ9cKIq6
a2MVC4LyPB4qjG0kk+AFXu+JvPEV9olRvSeJPrpZqKL/2wH7z4esQsS1Zt+eOCKFcFh9jrC79NfO
vHVGdwhyFScxB3E+QJLPwwkG3zdr3NGS3u3ZER6I+vh4D/hfP7Qan84P1kFLngUzHSkDCYzXWFo9
YzkMQVWEg1gzM/gJhz3ZWLsc/wObpGVeRgTCi4XUJNfHzOqL7C9Z45NvaXFdOupeBsgVJfbxgHDk
m4JKlrz2gSwXh7RdQ2DHeAOhTx/LqcIquzbxKlIJadkSWvZhDwsAsR/RrIIxd1YQTDUdPBfMrs3N
Qr2DWKJnMaaACEQHeObhXRvb+YLErm9OedJ+po4qlP2plL650JKrebqIxFynDd7baHummrNB6JZA
qvzHs6yC6JQPqL1PwDFOhoFgAn/MqRAx/L0n/5bRKyhFwf6KzhEWeBuxa7AjFX6TRj4lbF6qf5SY
1Ffg1r+qHugkKeNQtWfzp0MfBHO3c8Ut4qxJNN+KV8t3pRrBl7TL3jaOihtoupoTqXpRQ0BAgGNf
n5zx+Dq1tgAqSR+iFowH5TdseF19y7wPO9b3+QxZSegOEaxYSSW4ZmE2wazFlzx10k0Xq4n9TUfh
DZb4RbUu9v77GxcGyMYu9fjsYtOkpt2pNGzoGTUov7XLhO8Ibxc/7zNB2mmLhd6cpyUGSKifjc0h
jc/7Z1GUpqpsaYQOjGyBLPjUU73xTs0CqI6kWhAUqhSh/T0nWdI3don4Hn5FOFAe/CGNzehZ5aLV
8e4U0c7bEcNhTAji0J3uqA74051JxqoWr8D465yYB5HgK2ULxlCPJz/hrCmjetQIX+nU75UPxJFO
RLGcZC7Xd/jkQdmckIU0sILvFu5yoyrfSVNNE/h6Xvtxfr/gm61LYaqueKsEqE/ljmOFXET7YPTq
MJzHYkxAwPZl/sGKlJQLgAqYc5FXOvG9bIKV/5ZL+zEZNOOwxVmf4Nk6w+E/B2bZlogHEBrvVtyy
aGXhCXP+fI740LvwRyFiWCxpvMDQKL39PQ/+jcTCDU0dqxHqOYKOUSLvOm6EtaBRLiPlNTQE633S
LLaq5f6D+oY4SoRw5yBw/0CQmSq0P3d+1piVID9Ebp1f7iuI4HDmnAIgQixipLLsq79EDktL2+B/
tAZhggNuYxmDIvYYxhZ35R6Ykeyvtbyebpz/7Xzu/gVxBsRMkB9KkqYhue3OWHROCPK//C7cnpvd
ujLgTNdYs1CQCYxLDZPscgUKL9k8g1LgXnS5BCXAyGrJT1rnuqfSvynIngfjqNzHb1UWsEPBgo4W
JwXXkwRoRF+D+mE0BXnF2tTBYw35FY9BLgPyYBqCleKVE8ASt/06MJiF8e1osChBMnPJC3Uk6yhq
o2TCAWY+q8r7PTJ4ZyfhUqDYOaJZOwIGIoq2WJra74Mn98j12XfK3ZO/GrB2VhKvHgAftHUiNf2K
UUnkEcC7jFq/R/lF88RAPgOO6v6lsDyzSKYqwauH5InJsJ0nBUyyGmaEI7C0m2yvOqzBt9/4Zts6
KKMQz6PgJrwjQ4ojBrkAjVaICdW5vfIkDGC+ZvJqc+7yXbpXQvrrNDEvWHYWpvNRlhq9bBL0o1xQ
AGvLX9nwI0ZiTOBeqXsPXxwr7VzBCSwfxxQTJFlK3dyBgElb0M4yanpwM1kEATINIqeP+dzd8aqE
oBBDfQWbkE+aJ75hriBS6/tlSZIxmAeMvfa95D+V/i7n0HZz56H4tGOKWxO4Rm/ZfHL2AQJ9KNAk
C2TbdOWndHWHHrot4djIBUgtBvehUJKjsS+vsnjIw4YtylBwZ9Hdh6zTEi9jIe1EMiioVOB+SuJ8
0g7lQc4l+vq7adrH+UzwnU19rP1oPQN2ed4/G27rhi5bYCXXdAhj6QphnariGiDPc1JuR26CJlx7
8DPxJb17Fmda7+IlE+DDlUG9BXYtjx6xgwVp8kI9nIpITXRtqusesMry+9a2XbRUj82+tQ/G75vO
07NUagPQVHONG6Ysfc3Lf039s//x4Hy5iUeMiVQFNZ1uHFILakW1t3FKcMQxR7697QSG/Tnz93Af
QFpJOwZQQdfXzE9S4FXMvMnZ0szp7lQH8vVmJppqMicTWz48RENG21KitmwHO9I1Q+wFUkuSvQHt
mWbkdAJgYECFen5+HvPvXV0yQ+phd881wShCSZ+3qyNPU0aJSoQC4wL/LkhEPBGCfN939kxo2gd3
g9kdYLtlRsjJf/kuTd3rDUiDC5cdwPtS1Ws8XjWdKsJ5BLo8s4wqBewRLj5A7F1RaUAYTn6RxnOU
8JGnksqplWTbhqAHiyJXIcKWf8HDaAlT21KEFdz6uPszH+KpuQMcAfyC7Bo7uWOxZGpPmNMspamT
x/G1IlRkYQp9gshEnCof14uSaceJAXxZOJKGrOf0AlS6eSLI6LdFxORLTOPT47V/3FD0XOZ/B0mB
hygbAzKaNccfNy477yWJU12SC4k88Qp3I/TZ80SU9B+V3+W/hpViiOxl1AXdAO6RrI8EQ5UmCsaL
k7ntVeHREqli3wQo5Ibyk8fSgVNK0RW4aaSP/i6TJeiQCsUTmH0m6QGT97EkNtFkW+j15F7otfis
7KkI+w9uX2W/3QqzzmLMgJZPf5y1ZWkIgybAuvOo4kY0K37ByhgwvThI4NNcTrs2PhylfCRG7cUr
dqnv+5POdZorAdcNCoJLZZEjDfWYQs7sdalGlpPd1cPTtWOlAgtTV6kL2zjS/AlQetlhtH7uZrJ0
vS+FETCbdVYqA9eD9iYKIip+DsP476jqT345iQFj5XazOM7h+FBF1evyQhwrzABFaaijvIXawyqY
XvY2b0QbmzL6YQZZbGHPCG4Rhp3Sef2E+H1jpOyt45X8iszG+GaVGXOurzC3po6QIE65ir4+A+go
JJxO9RSyej3pjHV9VHYByEZC3FacruvKyewOQe6k+KmS86CWtvsXpdCO+JQHuLt7XoC6B7KsW6iX
ThlunVvQlC4ql+6xjoEZGedAlqmigm0+LcBzzdsO3qJtUtTLRwWN+JTckAS1GLP0BrFWMI9vTspF
Du+AYZHlPLpdCngQt4J/wiszjXL85TefCeC9rGRmI35SbxQJf/Hi4eZeFwsyrNhCI4HVmqUIlQ8u
K4cjraWkNfSll/PqmjPxguRy/3/wgGQ+be6DlEi3LWxBJusRG/OgyN6ZijVYBwxK2vXdoGzrEIm+
p/sf4m5vT8YV+5HrGLLq5ZrtSHlYjE0PElvP4Xec1LfmRF4isowGhL2LgVmHkxaPK5kOtz0yphsG
e2dRGP1LM/px1bwtuHnWn9FDW8b8RHHHAG8m6dqMVOv7mCS4EBzXycaMArmpydIIyV8G2Cay5v0W
jpdyuEBch+DBV8eggGwbfnwUT8gdyxd2JuZGzXEgTT+8V745i1KD+lxrEkOiQwSF2k/2VOWjSIYs
TQbbMFD6K081TSz1QWKoRulybXBp7STrTVngbaC43jToHkbqf5AF624YXkih8etZyFbbj9PGQvjE
Za4jjYPgBPocwXB9zhPaVg7XB1dd2OB/2zpjkgXl9mZ+sdQsESaxmvIa3Lkr+UoXVclE4vZvX8K1
ZrV0ORjB+Amj/BNixkBMkRdJf803RgxFQ/KQV5csoLNk11KU+vF8yo8OaS7/Zo/q1fQEfFLGGv9U
CRSr4RwvG0Wy5H4vQg2bBkkyrlY5frwyurUhrW0n6rf10+RepMh/VdEEFgqtV7VW+pZaQi+xYoBE
CStDqxjZuD5M7u1gcpRzDBvhyGg69oQzg9xhhws4lk248JoGJ6Kwtn0fMzMR7UJe3q/avRWA+Eia
VBrTMaAZvakuKWEU3lZJHHiJwGEakLEBrOxJ876D7QxEgCUMdBmy0R9gr1DpdcuCWJrX8RR3Knff
K5LaN1wZOxGtqUZsDD4rAsfztzg4pLhxZdKe2uWNHeSDy9fBAfJGUrRHhjBnZJKi7Nq9m8OqhgPP
U8CvTgwDJSX8WX/qxhXAQu+jYjdj/tPNo7v0Zxs2Vjca9qaWDpNsK0+dSip7aJc2evfmw675V5aU
XtztlFrsfWEfRDJr1FoUFoCfaHbDrs/fAclwBNW6bZCCnxRs94Nw0qU+Tnd5nhXbEEkYOzrCE/Bc
VbjEnRVLtGGKYHjVAWIkd6wJpq/rMDeH5TlQe02SJrwZXRPs3QTGkaP/xP3m6uwELrwTEk9BiVvy
pGO9yh/K4TpvdPRH0gP9sQmzlAKY3TzbxNGxfhaEO3OiqM3OOR4sTt/xsmUrD2tZJWiveS0zEZVV
RLXBvpSHugeyUqNoVAaIKcbuJXG8QV4Aow4wE4gOGGTd57gsqIh3j1HKWy2mST8lRiiN4hQetL4k
vV0xFXRF4Tw+Kmy3ECTJ359+yWyPYRCmdOVYVdKFihfmfj8PFONvRwakkVCD0Bdf/zW6NzdZuQvf
xSc33nV6Sq1bSLhavCO16uq8Hbm+E8iaecJmp1WXFVhqxr3UNXFxDS3PDBdjBJFyxkmogIdUmHkr
joBlCciFLjRgtzcghZG69w+Zu8wRv2+XEWcYyGUW5GzOth38OQgLAKy1Ue2En3/3umUREi18FIvJ
MDRthIP9FLpwKgy/JGBBFM0Fpwzhd9AngjoX7C3ZCBCQLcvJtRtwSPdqsHGayX2x7WSbhQROxBtt
IbL1qg1074yXl3WzrLtWG6muv63KQqRj2X/XXd81OkdmPPsf7z+QlTRl1kA9oPtxUm3Uv27ibFzp
xy7lhhzCvsif9tpd3JLTkR/uLFlH/ag6EGvm3w1Nx6Q9Ph5SFcgFgd8OQu6ABm2+t5KVZdM+R3v0
lqnqoWGcqFwRRqMfG9PdznQVt3o+z80FQDfZUEvUAHuoj1uJaueTHpHP8cWt2Pzb3YG+sB1xG5Pz
CDkGFyE6QMpMz8hdS7nYV0tKgliPLqHlkjiTfMCkVMyNp5RoB0jvuE6Jr7YYjdieo0BgweUz5/zv
j10XKbgmUKaX3y7bWxjWf7zojWRtbuuU4AScoevPBEr3OTX+NOPuUOl1OOgbkV6HTnfOd+XbGIWf
1EqZV7TEDUMeDTr0KGAzVWDWF6hT9mYwlCgyqCQvaiaLsrytO7gzgBSeV6ornp5xsTyVbY4Zj7tt
jjlfF5pmzTiappXbgnFBJEV61my9r3u+fnEwD0/HBmZvtqhZXbB0xn0AgRj8zWPx6I8VA2yu3Frx
EV00fUkbpVqMQLls+6UUvoMcbQAy+0XlQbCQ/3iZXcWNFALqfjpnB+dCqYFUBHdH/hTOITRKe/c7
XRQEhpxiwX5bQHXnNQPqGLt78hHkP8WQH+aWn+M5U3t6azIfnmmZOJRCJBfATQdXyN51lkaS3xGN
uLJEyskuS2TL3bfq1j+vMojkEFGdJonM7geN+VdSDN9dL6G+sz1o1UGo8KC42wJAdNW7N5efk6q2
jJTnSyRTskREv70Cne9vq2iEnuHxxVIuDgDk93NmcTXbb5yWLxqHjEjj2p1a7gqsoT6YQctz+FeO
Stgr7DAcJf6uNEL1EKSBOUy/Q0xGt7mgUj92XBZlyeSf1kGD9oUWZYlk+Sf6QUy/n4SzXV1paWG6
md2iQUNdfOgJ36dl0srLEoFYjTl7pPzTe3YcaH1U8eUWwAtqL6thOmEiqYxeuFyctC6qc6dwseSB
bMJF3q7/EisHKwQbP5iAtWjaVG/5Hn8b7D/91nommy+l2LC4swLMCBkhQWObu9ug7yVHtW+MoWyA
417zgyNehABC7NRjhce2JD77rNX6G8TcIajmGZOaXpXBslk6FBTAYziISldOiqx9X01y299RKQtq
cJ9wwomJSvtwfvFSHotaTXZkT/9fs7m+Y3ZdqXAmglg9fpyTWARdVN02SA3LjEL4K+2Qvkg9P6Ne
4hcJApHF4d5JAzmk7g4XzpQh271c0JTEykGCsX4WDWOO4eb/E7XiajbXsoorsCJQwOeOXJ9q18eW
Rdt+Wn630gMM1ReQEOG7cf+1SiUwfwzB4aGMBE/xnhUyF2U5JSnuNg2KcXAIrTcS8XlLk2LhXc3T
I2tzG2ck9NnzHJonjKl4OA+999ITAzjRbmEaXUsvvc+HjWZeLBDYGnKqn7MrnKwnn9Sijak+ZpBh
jAbFBSQ5kt5tbAqQyUMF8Nje0xMhmOORgRNRCwxOF0rFaHt30vsJ8RXVOnb/sgvcz+GeTrPBgOnn
PNTe5viho4QFgcebef7VV4mkyBEkC27mlKSXFGvQX739HBPoZCHJjRb7TdR7RGDxhhHvmE3RB4U/
FKg2ZzlAU5M8Vj65vaTwOIphzPydRxahjqfVB0ysAEl2fOMYDxCdeBmF65RDtkEn+oGyCDIlBq1x
I/Kw1KurWvsmWMRHovMMp8QDqUICfX1SJduPbmk/IdXQycsyJ2e9tRDvp0zfiWBjpUZxIfYAZcTs
DVLdEmfa6qJvXdY9I19z05+uNimZR35VlrQCGhXVAMfWRtLtPbK9h/5adwRdq4oMQwumP9UwIsIH
Zy28kckIt9uQVOx5JAgnQLSOjCKz8ihBpIWBwCC7jVQNO6qtApYPHjAo/DDiogkmqLuYTbOFaPo4
TCjvgr4HDQWtAccRgvKjw6e3o0YHjDm/jJuMvouaHSiApH2Oj85ebtC4pYjWV3bfkNfJAMDR5dP+
MXpeI5MOtbvg2gt6dzXpYxJ3jr7fn1CkR4n2q9lAcgB1iY61rnvWIXkbWsz50MzCgwhou3qIDOCy
DNWT3uRuIvUIpnZ1iSSwaC6yRBlPiaIeKNkNjyPw+Dwmj2B9Ipct26EWmKh6eVsO8u8dBHNBgkgK
QoBSWw9t9flytrk67OMcr1RoSww4Tsh/85JiVir/FCQ4vjxg2oL70ctNjW92kya1wFZSlssOQIrf
wpgiySNx05Q9DtrcyNLxHoye/rXdApC0iKBmq/MHdLJZ7EY3P3xJMK42IiDr/3Vv1qYnvw4+V0MB
lQgPbEo9gFak9JxI3SP+fNsDGSkA/fjc0AQ1axBVJeDcljH1DISdonNyUbK+zcIJebrRnxFN5V+f
3srX510o2tvK5Ob+6uO3YKeINA6bi1vEgHPlUWmMwoakZQ75KpSr6/byqc7b9pl51MBcJfCFE7QY
ibnniNCD6WkI6LRq+ddOAwgQ8tmAnJUAsrJJA0i3oHoR+HIf/4qe/y8Ad9tF7lrCYb9S1wLhV1ow
x91eqYvYdkHhP2REQ6I/ls+rnkGrZDrzhAOHa0g7BZaWyTY3nnVJPiwVx8H9q7OjlaNj0gRb7F5j
YXWGjSraNMwKl26ukrT/Vbs67Kp6OW6NYMsp+VIrc+0W167nL12Fae68+gBwzmW89mXuzYOw9PXS
+vQ3LHN+qJqGl6ROxGjyyhRfthKTSe922Z2lkWnFCNDzgmcbAZNFY+o0LGYp4Mf55vfiB2rP/oPi
krwokb5QWlH+fmXqOHa/xQPIB1VXYbwLx1xlUlXk2hXCZ2ZCCmOsd+4yc1roJo8GeBp6zfxDe10/
RuGwFRIifO32KMtWXD9DLv5Y+NlRJN/Os4JHAsok6y4k222aJAEcymgeRz6SvU2F1rG1okCJxE3W
ZrThrhSOMkYV/f/TqhJzMiQwfdDlKaevG+roLLoArJzXN/YNCRyjaC9fMGydzGVmip868NQrAGt5
qmf2FA/DwqdQNoVkRXhG0RXO69SqKc4QLEGSObpm0PIRviqUMMiRhmdg1UqCSHC2mPy5ypZMRKx0
NFvkvaUqwvEs6BHJnJHgJpT3O8AOSK8FA7sj/kHfIMP9aKaNhtEXZ76iNbD315v7oZQunCpzln1S
G8DAuU0adReNFlWzcom6PnT472fp2XheEixQOp6RavMK4E1W06qBOLOEFqMv0poHNCF8phztOg+F
0TqUMiIGCDF4D+RNJzAytHCubWlgLnkZDtTJAo+idUP7jublyEHbILz7X0voW7/jGLLH19S66JMX
AELmUo0nUlgPb+wTqv/P+dMKBMPQbMlcH/o21iuA/cq+2ImZgHSM291BaZL97oVoHxsVq1yMYPRJ
xi7EpoRdhlOTVt7Vj4O2qj66jLDkdPz5GrOoEWUGRFZst90NMYrc5Loaa40pHjRCzwQ4lODrZbiS
DpENaOXUeYrqNUeH0eMvM05WPY0sN+Nw+P4ueZUqSiNYJ+m1dOzz72Vl95F9M2+indRTJ557d5/P
NmeYT2MlekVR8gnzBrYvitRJ/pqInfSIShMDW5WjcPpPlUhmIXHCstdwVA3QwNqhZIbublg9KINw
iB61jjwn4IivMRG9e6oApt2LA1ubBIZmQDiaG9sMBNPlA7vWyYWu3pnQP2aNY3TLNXsSYi2OBWe7
rDqnqj4AhJDRf+aUTw6wSUWgkt62PGd9Ni/dfDzNTVG3b8T/Doq9NZjv5hhutVwdJZI/Z9xBIyqf
gr3zfs7r2wsUkhnt0mGvKmJ+imFwA3p4i3yLCuOYZi+fLKF6lFGAOciPasQGykSNBeEBH/Qtad7J
ZFhTjzzZAvKxoHs2cLw8FlHOf6+hrBqxZARl0yt+fkBkREAGCQdznJaKPJ9eKQyNqPh0LmLDG+OJ
9ZkgAo+RzEpeHex8eJD781sRIleMY6/42pU0xwUKdC2CFwpsgMLhqk22S6kdRoCPhJjqxMuE/RzE
93hMdcsBgvy5Tar1i/jup3XHCwazefEpR5PAXGxBRv3yy6lJ1+0v3k0xEgwDYMTcTwIEOw6E0pkA
oiIA1yQH69yYuQoFYHQ7kifam8lWWsQ2qhXtCW5oRzXRFvrkpKB7OL/RacSneaDBJuqzPXB43Ele
S9zdgxbDoP3vZtsl+sa8jzhwCYuDxSO+VbZmn2+xw+MW6S6KsB2LyohvfD/bYZa2K8MyKWBxOiaX
9T4wQuGbGG2wWuHy/eRgAoToIg3Uj8Day6LDITn52DShbj5BnNTfi5BmGZQ9M/ZNDRVfl6ELkp7/
ZCsVMlPtd+hle+F9fdZlX+fUcqdwAPt0R5RgtYnYNMIkumgXkl5o90PymqTQ7sLrDLbgHXEuUTiY
UIQV49nS9aBTzTlCkl6a3kPZFUZoYGWPAT1TZeOniUQJMnMg0Un5HmLkhl9RAKSX5dZumf4sp08g
5ps8sZToi91HigqP1GwIPl/X7FUzRBaz/W4bRKSYFsucRrk4gpjtecjwYz885LN++cn+p40i3Cm+
B0tMJic9BV6ZoPs+uX3hCguxl5qlpKU68Ye47jDUFHBMkWQrsA/ZXd7ZtMt3iZhhS06/zYVqJdW+
r19TBJmEtlwrmQcWCb3DXi/+M4JNMsfQJyBuI495+I/3Yqz2YLkBPOm2lpAPj7pV0mzZ77KSMgt9
sQhjaTd7Agk7ILTMltonMHRLvAt7++0Q9MTlSByLPHd8tiEZpahhjpKpE0ZQqGOriePVQUCoT+r6
VcaWVmZ+7SAQEThfKnLtC24VMgK7MEA9DenUmBtc8MpFIiaaGvJ5xSiLuO5ElaGIHuE9N+QU2NV+
/DcT6iiy+bcrp23Zn9yCeLMFsXCazQx6XrIb+93Ei60dT+U7MJ4uFFRQucCg0o+oTNuvzXmE7q56
N7ngfQGAbuUmBCz7IrMby7eKPyd/5aUHomvwubg5v106tbzKU8huJRMWuuSLdR/RHc0rhA4S56J2
BD9UH9tbMVl+zDDLEh1Ti2lLCQ5FUVb+1PZYdxTRJHCrCONGq4sfStDO97msJ9amLpJ+on/VaZKx
GFPcVqAkh8DDNLuvF4j5oeKE06YY7GfW1nS2pCVNcxBK3EtPNgNuWydvAMOzHJsF10i773XoerJz
ViFu030uBPEMrt8YlE48u24UFukQaIAZb0k35fHKj3rjxpicryFF9Rzf86rmNeWqFSDMTnhT8mEo
8C84SaFSy5f6IQTMZPxQysLKeuC4lDrW4dq9TsXcQ79ceLTwtkAfjx4u490VYgCzFPz16zIX36eQ
yD38rWp02sekw3pxY1dPzbhRXfeC/SWWhY25P/r3EPHgLcr7C7cjlv2PmBIjUcnh6t+tk0xo1j/T
T097EsNJffDNd87TAedEV9T9+bWXi5Z5rgewjP9RdIB6wzMa8QnMGcBj7GG39JqK1rqWyqCMPP1a
/ALFdFFoHoe5WyAdIUB7rasby2pmjdaiAw9UrA2uNEhCrmzsp7EqqNF3QYrmwbjnZW0MGud2X795
/nX64Nrhd5tn3KpIHWdT5FGM8gpL8S5+yYAAndYGU5el0XRgPianDjBfXt9NWDI1rketBOmwQAVf
FrFlxywGq/Z11UmW17PAt1QfBq0M5NljFvsn8VD3kMtQyasJOqIDLRa3hJOUBPepLeCVR5wIJmJR
xz6YHTWLLZ76vGt4Zl6d97N2vBBQrHVrAgTLk9ZfsaU51PXBSD83MFF7T7+64j8WZu2F6eStsYH0
bq2ddQ40AnQOcx8xbSWrVspUC+0RJzlCANT4hfg07J7tCc2LpD1+tvLO5J3Fjs2h/wBr5wjvoaVi
K/adGhucnl1VmKv2w/gpJJVZiorxAzRx0TgFu05pFpoFAZY8YIbOSWxfEnP8lynA224kEgM5Rs8P
jxO9UY4euHSImBhmolEhtzTkEwynluFRVbTtmHQJ4urRDF1YIdFNLKI4f7pspuxJdV6xR7K1XO4u
WJcluoxJklgZNmijNa85jPBxtqpvN+IqBCJhG4Rks8u2HHsglYXspRpZeBLppiWICdDkUlH2S1jP
QYDUwGHuBhiEM9BFb08AmS55XzpLDeP8nvhm7X95+brYHJLnd0D0dfJAWp3f3nQIkFN3uiqPHRrr
yjRZsLq7HYGwP0bqVOo8ianaLUJC8/tNl43NZYbhhCqxdAllz1wb+P7X3sYKtWvQGAeKlbH3bgBv
Y4qmP3q0IRE8l9qyGGfputOBXcdx2M+iUW8LhpYd5/LlZPgAPouxZGR88CAo85icc0xm2+J3VhoF
CZ1nylRbVwy8mDsuWcTpTqGfNQfmprhk/XLajhdURUNTA5bFpn6Nrnuu1ADt3/m7CeyPeXYtM+CL
gRz9A3uOnzHnIqAIocyj34/SJu7o8y06LwlnH9EZu4bkUMeYSDrNEn3LvA05mU6derJ7WFQgW7R5
TU4bWmKVzDp2BBugkLZJonwGEX9x9GUSDCmFTL5NcKu3YyDEHciPY8ZjGr5t+HKPV6dqaJfW3IPu
Cnh/n2u1z25yPt80A6Gw1f/Nzn2kRYjcedgkPM8XXJmzCXQ9HahOqkaJ+E7mrBpaQDHb4wOOONtl
iK+nLz+2xLu0RnO/xg1pxLao/cIFKcTV1FM62vkIF3X/A3Tx8oujGGyNhOq6dFjY3quJxFZJ5mit
UfVzTz3TupuPbTZoT/6CLbGm+mcMxwDZcKfJMqqsn1l+QRQNeSh9d5o/cOSB2hPwjkw+38pYdD1Z
7Zvo9gD4vwPjUfjsqiwVbNXQGGVrv9Ie4O/mbGMkIbVQn6pYCgovXPTp+p0dSOx1YHFUnjKtZfw0
emuY6b6G2OkMWKlvYYaUh5VabfT/njPI8qdGSX1o04OYxYMc7bljb2qP5EPZakRhUh3U/zWTBFam
YkVMy5L2/Ru4EqHpca5jF2N9zT6iwl09a1wwrDokpYK1AdkkTQg291qTtDRw+vrSyYOYZcbg8Sqa
2jYAAMJ9W0B9tp0ajMPDhDUQzXA9gHP273JejdL3dD2Wc5dVbFIrJldc/Y5bnSkznMI/Go+LBUQn
7EUT9bnUgVGSUM3iK/FHOgUH/7o9Awulow7Aj0mNecYYGKVieI8II+6oklZu4JKSWQj4VqsUAkHT
LDksapeDYLZ9nKW0bAgjysHWOCFINOnSwcnd2tocnz4cw0pgTVrrn36vygPfsnSh6v1sdIGViQkQ
2bRvwBARiVwqmTpnX8FB7uPI/KHAgHNypsdsxW+MB3KOki5xoAfjweZXI/6KOyHj3cDzNA+yot5a
dC3/nKUvUxY1k72uxwj9myqbuL4mDrYz6s8sicmiXoXyOG5ZSS40VL6FmpuDqg8vU/XOc/3ECG5r
qjoypvZhZ/b4u1SNjDfuUC8EQHk7TJjSli9aNCqBCz8V+GhzLF4M1zvCWqQ1LKiZYQRyJrZ41/Vf
vPRKBib3+aZC8HGvNzNG1YqKKyjpEOsRhS4lHAWNDZaWiRvXSIxlTtKLeGUIlAFKOmVv8Wnrx01+
uvCQC/rYmeBFB/Yvtc4t+FVl8ZiWVuRYFMf1tn15hjZo/ho696OGveG+QPVf3Trv2IFyH2Y3iJOk
uWyldaeNlSu/L+4KCooVgeGTSquWEResSOl9akZtRK576k7v1y1VZjGH5kKTnLpQkzjyo0uiKIzy
Efp4qFV46aldjDuWLI/bJuMs9yxdkgDYayzefBK3PZnZbl3/AY9lxLCUVWHXehp1/pE7RrBPrh+q
PbA0GnH24EeKgbzGcmkujlNSAc3sEwK9BIJjTkCThk0+UDDd+Q+XZikvTjgx/Dy3R34Uly+OCI0i
Pmqbv5GNXwNnB+OzgFKkJ8oD6JeBx+AkhiZTPtylRkwksL/ak6aQJvUkCp72MtPIYgOHVqM2z0Ee
Rz3PKVtYnCwhxlU41zWLcz6TW6owcH0nTOTzaMkO0M2+TpfD6p7aiqt2NE2yyIaiTzCS+0jOJvd0
VTd+rFtkRK2mkCtrONiSFzFcVLvs5yZSJ0to50bCbVJXjjNoQpMHhhWkOz0T2WhvyMpIm8izflrD
pYs0Acexg34txdepuapKQKweSL4pBoZqRkSVRBkQrOQof5+5EmlLHZ8msrJumncdZZOTF98qy8lp
ostsZSaAi9EwYTR0+HmVY+abQUhBq8XP1mAKDrt1v2MSZCylCVDV2BmFvgfbFc1nMpYn3+Go2dsD
NbTzh+5vL/rpjBMDwmUkWS3qnGfK1ATDw2mCs933OyxCKz/jmKJvuSkThD1NwfF0h4xmCyeoXB5j
zVHKbokAatfSUBVBvb6Jwz9w1R4Shk1UXtOAvC3vlTZQH2kuZvrHLxd2w+Lx+Y/RPt59eXv9jyYH
vJ51oYUWJ3nQjrALsLoxbB1pdsVBR12sPsPLIhk1zHv2uPzmXCgZMeGiVJEmMGQ5Nbk2ZPfOmcBL
menD8YhewpFm7aJNx466Ol4FKpzCHucnDKYx13/+QE2uBiVUrcHWf9IxxZiIRgdObjpp+vPFLJNT
dp6mkScegeG9QkR9rIqWWXpEznmQ/rR28AbMX+NdZLwx1aasfiuFZmgxFuIDsfKzIC3eM5bY4fbs
aOgKEkMFj7eIrp0/LWDVsjuC7zxHRbaHjSi08uyKOgdGZIYOwAm1roGMXu53Mg0tLNppHNd5vaQN
ASM2hwOYUafmExCTT/P3zYRJU46bMyBYuT0qp3yLh77PLS9bVBxlu89Lf3501dsrgvJT+K3KoL7A
6idCyfr/ewHAgwzD5yeSyU4LUiRvVlT2SWzoJD7v5J62jbR2JhMWTrAxymSZwJyfs5lFG4WC4M1f
39mjBpWt5DYp17j6MptfdUG2CJmdjDi1xrrhCIH9QFvgSIk7Yg3mqUdx2uD3Xwt1AYTZJSAF9qsu
UBspbn9SJw8JA+19kWwC2uX6pqTbQrzP+njL2kQsxlMtcmJIlSYsXON77CyB6d81GiFqeLdbiSJs
eEO84GmvDNy75fAFlBUPLnVJUj0uYQPeId2h0ybKAJlaCI0tde8dCpZIYoNoTvYw1byYdh91dqyU
Sy8miZz2UNizPN7Eq3RWDNTYwciyNybJhdlqDf3sp0e9NlzXhKzFZSjYMPC2iPmzwkLT+9ZSWaDR
8ZFk0P0vAxMZpy+y4WqwmYvGUlHA2muLFOUh3cQcoMWXGOSesq8o+B9JA9UnSOPQy55LE0NFlGNK
TxUyReGSquAkeamXwjRwYU0fgOk2eR+skA7pZ2Q/bjxFpYtta7IGASuIcz52Cw50/3lxTC69CWcp
4VEYB4xIPIkA0v+n5UOCpJX5y0a9nXzOomzGepChsmt6jycxfmUHc05+6m1zcnAMuegUsfykbC0p
cWnSIpVf6U82JJl5tbn2r+TOsxE9+9NVQBRiaOHZGoljlTO+79OumQQ1jY4TYfKBzItWhbMPVzN2
y1xf1i0qXLgFZx8ndQC6vpxJuPI4H6YpsGkKayvd1WlZmYAdswge6TXadcOfSnl3hRKRr2YELNUZ
2wyCQRHZK4D/atbMPkikxmF4C92xh64EVj7+QRz9VBMcOTXZb4GmqbDdiUCj8jST9rt8Tas4cdBM
gcEyy4mSGoZzoWxiW5ma77EoSg1ey/Cp31hHqh4WqBqj6rCseJa3OB1m4I2d+mXDkW7x2PCyfDWc
jAiDcHrGfdC5Xw1IWMsYt0nXRo3WR8hkQjXsS9nQ64cB5DWNFLQm1qcD0Yxwg2k/MX3vuldGDNt/
SmKPFDOkt4U/YeB/Q0JvyFu79Vq+LPanFVNby2+bSFWDDM4zbH06OZ1dN8IKdg8A89o7BQu4VqJs
KjUCIVRBGYbiqUNcWIWL4g3Y/WkaTjoyGjhL/Yu80Z6fZbslV6EKDzXdF0L+p41hHrzsIyvRxTBj
YN9U3w9MGP0QvJyQYRMaGMgMSUK4D/YQAYbziRu3ppf262wtDwUFyJ9F3/Abc4z0PTFIz/XFkgP5
lgQW/yhYCa4uxNY8w0x4KpvTMs9eIGQXLKseYu+qihpXzvL9Pq+hY7br08nmcqK/+blQjDCxGhZ4
cmSUOr1zMvDBjE+8slrRGJpqi7jTvkbLW8fmLTQG6qJ0fIUz22CjBJ4XLmcezFrH0u0C22Kz8uxm
4Jxit1r6Gne5NRrAsklBN3tYKdeFcNQLZf7Uco7iZdwkVuxJUkQFh3ipyMBIJsMlFvoKcykAWe0v
TS7WrNUSeDG38i8hs2pFLoRGiGrmdo13hLCDotYyL5pBnpYN1Ts9Ic0w5CxP2jGnm0aXDprPHDdz
L9sB1f/NWyVuE0jIulJxBMGgCpbk5EjCClT03+Dp/Pzk9JJnZIyJPqbBflSq0crQUMt17jMfQHYr
5+rcgbNHY95nv2NfAx9gkNNorBOAQKrHM6Alr/XldNUl72ewj/eYptJQtLx2YUUU7UNa+NoQ3O1C
Lbhj+HeYYzCP+KtPTehXY28DdPLN4Ozai+h4rsmHS4glONuJ1oATAJ+m8VaZx2YgSUzOoNqKzVbN
wh2tJE3a46WkU85CEPi0ZVXvPtuJRTILrlSIwHXes0Lt6O+PwRdluwwMnUw1da7Ko8YlEqE7CFL0
5h+UQnokQ0ZHL8EbQTPvxK/MGYkKrbkj6A/N8jKF9Bgc08F+lB7Z8OGDqDQiai/CntNZOZoe9FHe
//riV6YUuoni41rgzOQc/KD+eik2PvhcDBuuqAdIijw7EUbh+nTueBVMsZFQKZv/HAOvJ7zl8mN7
jSTaet11FV+GNPEO28ZtW3fl5kShM8cVsgReYYlI8yBYzMPzLiaoYEE0PdOLz6XqCHNzr6NEYDxU
f6uSztvaw9c3qmiA0SRrvqc602+PE3UBLtN5qZXKe34JqxAlysrv0MiUg86Do4CYiyDGrejuFRps
e+bEgM/LC7kdd3K1tTgHcPr3MzCCrGC65SkchQiEEVhDhcNgo0ft+v2K6Et1w81xwKgvQ+9X4MPZ
h/k5zWAlOhMreqzZLHbnS1mYD+XL/Z9Cwasgmq3BNLC9a3RkNe4AmeRwwXTPVHQWNx8PyWftJ58B
3ythyaQJmqdYsajpXD6RLQQrhj4YrRuu1a36DruN5Y0GGUG/JTw8pXb3JG/gsXcMHQ2WCFN9FOR3
cvlFvPLJXYDccRK3fGnvAxkxIt6ciRPcgfJ9zYmdW5W7MGnvBtqsc52JUymptN4wJ7tPpGxTGkgK
GrNgexAcsIofYp1jMyOW8ex1usHh1wQ5jq1AMFT6syTKFcICbqJEU9PhM8fTaZtybamaLdiGI1HR
QEL+RRJPIvXY2DFRbvrWzXZ+Pb1+rzGMJJNIgK9ZOld26gT5EnJ3q2g0n28EdueX1S9ZseXpuYhK
BdDxbEEG/GspvSsjNp5wNdgDDoiOhy2abN7k+RTROnCg7KlQU/1SOkXkjvQ0baEXeq0VQztoOMxY
vM1X6QncmfDV0AstEoUtbNUaibOW/ZaGzVgohLvfYhSEJAX6agoi2u4B/z0IfLpwwuKW87nmBPdK
Asa+6okhksiEUxT9OQI+TCcnwRV1NVa0uachOzXF+mmrLxAW3n7Ik49kCDj2a69NqfrVHo2fGWTX
rEGsuIGaYL6TCmOgJpjPBG5Qd326SHGXnwNxMNBMkLxSQWDOj6Vo2KhXdRy+bLzP3xcm3J5xjSze
tCRZ/+UQy1d/gcRG3QyMACZdzEOx35DYVGems+Hq7qZ9xuX7ikuTAtdqzFFRAy/d7MXJ3v/Uu2Hi
Dtmyn8KihK9rguN5kEJLB6lu+YzXyKriJegYFbM3OgQnoCNLy6xjDS0c4Wsdk6YUx43NCP/4kFv4
NSIP32N6kfbB43MocsZjMTdkMjaKoJbbuiypjfG5yNmwcgsZwp3SaCgUC0p5k64KlFX2BmuyMjkI
HAdmehGmEXiBEyP9PZpR2StbmfNCxisz9WWeGeuvZznGYe1q1DsryoAMSiwRMT8fTW3H9Sya081U
9ZNvpnTnRQOxLJm9kzddCPExlYr+Htx7QhKzVA2AHmOQrGcRiyv5CDZh3PgQaKFSbeDlGBC5diWn
89G2zlLvQFq8jkJe/9JIliFf0KZFfg4Y1Halqt/SZZfsREcURdAez5wLL6G7ZrVK1jUQ7M66NDJP
aMmnrOYahbgpFDCOOyQ6S5o7aklfm8/mDETWd41JWkL29nFetPZT4wC4QGkxXfsrJVFeD/PpVKpF
n2zk6GdAiddpv/8shrPlp98+By1RXEgLgiGqcqE2tUMW+9pY1o0D1dDLTF4SBUbjcAJbwRjcAQui
FbY0AAsZFWMld/wM2ingPVItGge2ztd3GrkqV+z+nMoA6FRPvnLpBRJftxGVeXOWo+djQCmSArme
DwZ2xlRXoiNxEMcMXTdkNJM4Wkw9jJMZ/O4QluUeJ08Z6YY2TRK3Ek8YnMxnhbaJbdtwPET33wzz
sVLWMgK1gZnYhylH2xN2QPyqgJskq5L1LtpmdUsv0ueEG06rQzk5zXkXqHYZZ0msVexjgjTrTuKF
mFTaXzS2YIlrvAZOHGUJ2wC2JfE6s2qxkfvxMrlQBfBZn6dqnpR53qSxlbsFHPFQckivqHts4KnU
uR68EI45vOtYwV5UzeVumwZidTY0z0sUMzVXtBWe/oqwY/8Nvu0zU8tHBFvx1twyXtc+Iif5yzNh
jpr66yVtMZz4rHZ14E0aKiWjAdvKd24PEZQLxcl8do7Pdw1ioSbOY1ZX0BZUKiQNPLBGdLX5vPMF
URBBXRcxrFQok3fdKeLS1CfSvlpTJVmalwnCJqLSB/S3An55RIZ0IiBzcGNStMPrOM0I2Qhci1q9
2lis+YmKQo4AAxv01AtiV58OoJ6RQYRuQbiSm0EBJOF8mHiTqXO6XvZabUlOb2TR1DmAV5/Td8m4
t26y5z3bN4oqs9cFIzdEVYHf+/mqPfeqtyne/zgKsgyuVyFMECBgjqRWumA97gcZxQD8ilJO6ZMH
ZwRU6GSUVgqLFbxNK+fu297uYvVn0ToWivdF/T3hnTkwjRyOqErlOD/adlDml7uSRxfNpaNrRmUj
rJHkLZ4ZJY4pQFx2Yp2jbCdfBDm4hLrq/5gZKKzqwiRrMoBKKl0QeJ6ZKYUy6QyUw46juzomSACR
UPiY6ZmsuDfWROvKVIYhfiAaF7lgDVhjibTW+aWn+Zykjuz105TfAamguZHb4+txudat64+sREml
Ucbb3QrahIPZmHQGLCS/ItOzfn9BJz6iFQGnbFMLiZMb8y0i2ET+Q/KQdF/ntZt0UEJfMBTKtNrF
XMkwa4bNh1Aa8xaYd96pP1EkT3EGqZj2oQnPnJFw0hXLkzbKSJNXFn1us3h9e1hgLRjxXBs4Uciy
l7rVDQxPNPrtxIepByt/10zmwMOqJQbWcy3hOvLgwYt5kYPsJ3wXS7SVsnys8yJclJWRgla3+dPU
UGkdm3CC+ZSWHVG0rD0et2yECYup/m51CBhxDQ06fGiHgiOZzmcjp9mQKM3wKwaJu+PW3Nv6tFTE
aaH+ctv2ag3IR+obAvOI8293danAO0UQyZFNzVS/89s1zv/fESLFSNKx0zu5A177AdMWotfAfzzW
EvYINs7lQRiSWXk0Ne8D/NkpcsnAEsekv5OgBlPKUqZTeEXhAOLPfcfU6aRDhzjIwjOM+5nDlcI1
6xJTMnWxF16kJZDxh2Fbzs5sQXDE1HOpi4UCdIKmy7DMU56SsyDtmSDJX0szzc5xdZJCbOKcXvnq
TgC6AHUcNDJMsEjfqcMmXkNlRAhLq5BkXxfAFP8yjfNXeSmNf0GaWUTXF9R3Ltptou6IAb1qF8F2
lTO+QKn487Tj6vPCr6yXLyolVmXSu4IEVcehkpowhFUmvLxxneXZr8zY4lK9BWMvKpiqILSu3b2q
GlPaNCqW2/C0Rlo0Ery0WkcZRn8i0PWOdNPT7A3tC0iKY3F6peWDMKKgK9zMTjRhZISK+26YuRpp
lrmujDBda7i1RoDj4NMbaCxTJRgNFWXj6G4+C6Frge+Aytla8hlNqFEK2NTnTbCy08bWlEdZ5KT0
NNVE3KOYdWj1Qiml2npU7u9eYO4E2b/aJYcKN18cg3bJ459HY2+4DOoP3m0veuwpX+t/WeiNO2cr
i++nokaqvrrMtVCPBL+GsqM8ieE+GNBwyRXWMdRhT7APSJDzeXr8Y019d3q7ILyZ258rTm17qSRi
gAbZKwDTMucqRiYucbkwIMdv4qwUX/c9qaLH6xG6hDF0Iy1cBiD5DL271dEDFlLyaKVI4+Bhi5Sb
uyTU9cis52sHY9EtRTiSw4X4u2trV8jO9g7lBHPOiyLGX1Xk2Bs0RkF/jlM+1M01FUEtXe3vhRAd
uK6ZSIPH/92LfIQxQqJh7pubHeQKNcFengQujlTixkpQ9OrwRNgc3uMvVcLilglBNWcZlhCqMd7t
eGnT2L8LKF0D6jVSP/4YHTKB1aeADQyB12XpAHbIZFqEjbcagvi8NmjXU0eQq3kV2OoSw6zr4kSJ
+qZ4PiEJWpk+DYSclaFunIAC96XVdIo1as9bv8r/FaSrC8pdS4dZQeFgU+2oKvm8O9POXVH4WXNU
OaRtm7tqqAup9detWW6x6dORWXZzd/eq1qZX+GI6XY62TRsw1/v+ljx6WqW3xIhDGkARio2FVoFR
u+9tQEy32bIzKp1+qCEf0hajRlpcOSrvHCZomUiEJPy8zD3d4cD2QV10HaKm3ObjFfYmPW9PgYuO
2k4APZ2PSgUo3D9/Ys+ANTKysjUwNmk9+z1bjx0IM234fDCgRfqON4I5J0VS5QPCAxrqxtimISe5
dQBrl+YD4QRyupCnXjiHG6xTunEJVma+oiUwBaEzBB/RgoaDsKKhwPfVU2YhTfulwJ+5MZAoUopl
NdMLYKk9bXudFF9ikOGDOWmS6WDRRB73JC6yBd6FXsEFDxlBhCsvkp7MqyR04NEQo4pzOtby6Vkq
IyJ6fqW0uqy2pEnnJ6Mksn0Zy8D+nPsnc7YUl1H0WxpVXbSxOpZgVObw2Ipw243cLR5WD5n3BlaE
odHAf5FPm/8rN0mX8Iw6IAkZRHIY61o3utEivgcrXeTMVfRxk5qHFKwt4G9c/DPsNaFgWdLt+Ajw
SO2g67nzmxQP/CYZQTVh5u0NhSkijOQX8k3S11sfoI90YkFkrRDK+H1FkAsiuhrELKKQ7aSXR9vW
QtWZvzSIwSlXup6qleafGikgDRD6qZIEJQuLybEBV5JQNYvmIu+OVtbN6UZ2Pa5bHx/uXOI9AiF3
t7pU3MH+dbMsXNGeN4uIfn1GwV1BiZ5W8HI62keb3YZkbGEU9WIQwKxfbhnzUfLsFNo0ofLK2Rx+
TAX59K+I1O12CpVTx3kmzICZ8Jev5hvbVcpan11D6DSg/SdOXW/3NRZG/ppM13HPC+j16dT2juy9
VVIr3Oupg81+bzCuoClkWiCCVtTwuAEz+vAXHRZuhqpQpbruFjqGboPPGqF/dBeIjR6kygwrFlcu
Urj1+bJil3BThDyEIUnTRBH+b2A0mrwVDuX/Ohzn9qXbf7f6Q44NHpK65HeHJHlMuEgSOJ80fItC
IaDmbW4M1sFtNQ5n3UM2VmqhlXc5MwGUj6ZM++auZRSv6w8vKYIoePmWd6cZw/5POrNF/tw75veE
GVzPGySCm1363j+VqhJULeVZKVfEKpyfGHuSFqMYoY4IDr0iz3P6fz53q0CFEccMvS48zZaKrIkn
8c7FtqsDFa+DiwSZzIQPWC3z4LGoTlMAPYx2dWDJOnlB/7NSp7wJhobH3uFRYTV49RpOtbhicPcy
DlLhxmRMBml94ATVPRPPcjKT4OtKFQ8X3VNWLD0fjnMtHB1VwuVIo0/xsTZY3aWUVMGUtU1qAw02
dodD9fp/ID8QdHBVJaNrFu7l17FDEG1IZaGP8W9p6kSUncp20okqW3jh3ilaRhTHfOQAvX9uHja6
sWwqbtepPZYNSDy7ZozeNerC1bymkRmKzQl3n/8UdUR+jFBKzwIXa4I5yKJAUspPz1Unf6UMbNwf
SKOU/4MyuLipmB7elnB9nWjVD9sGhleOAz6r9z1tbj6/nb92MWmlJDy7aDm6hMnrNjZfMARRjqdF
B+ZdV8InMckQ9mF1t9heOeDMSBSzFg3R5ykCemgTVG5znUW1b45P2S//C0O4cliqgJbapyesiFPX
k7w7/hGzRMByerXq6ryXP37rwE8vKRUCZXyVGrjdtHfVWlaEfea4cFdzrNScQkC2aUYQwAFGLAYI
ULaOVzO4nC5wa6Aiw/UsZ+haWpu6bXapkqskUiJzVzbcRDT1qPHmBGhTrAzqClhrigIPHO5mVMHo
VSZ9ddDiWnYyl0m2XFHKxDMDlC5V2si/njPw0az7d40PSFNblcEaYRHaSYzwaRFwBAohco/C5/YM
SayVJdUAM0QvPC8ZOilX7yHe5K0ZfXH3gstqIxyAD2bzXviR5FbgnG66qFGTAyYSVlzfdZNIyA6k
Gl2VGi8tzY3zkz/82TlT6nbQ4qqXx4LtmLQgZsGUIK2DuajitCRhFuuF3xOcv0XkDDy+6RY3d0+w
dhZCCzd0LIbpXyXs4u3dL7Vc16VD1MEc5lhJW4t6LTAFwQiabu5n90dcrlTq4UXwJo/vPuGiTo2+
2PnG+exAZnCo0ao7Q40vDdJY2q7++a1c+49sLjb6rztyFV8Ku+KmHliWUZJ5SzIAvbaDAX/pOB38
Awppn45I6GNEW3mMa3rRqZc6bN4uSkTkQlgypezd9Kbfdr6b0hxDI/Alk+c+d8guDPQu2ofdqgsh
GgwNA+4/Ll8nTn3ArQuG81ggDz0nzdNbwJwlmzOsedxDyRTw9bcwhWPqPlk4Dq0Fnf3iMvgmcS7z
Z2A/pr47NfRclw7HNlE/cWxbKVVRnv9Wxu482Fd7bI0JEgXXpI81oDzY3WJfbBZbeJpIv/Us6crH
l6Z7G6Qil160ApYnEfJKLxyKI6NPYNd/xAPaGdks3dpxros9Jw5ZLvXk1eT3VQHOwaapzPC8Qdqf
gMDDmOsu/tfplaybOxwPIS4xeGewkse8/QcnO+EDHHtSn3qJKrpommDz8+mIOVSpUcp8efwqnLbN
wksrGRYenrPbYRDvHng9+vU+bdTuoXo8DuE1lLmTamn+Gn2JPvMrra+lEnuborXetCzKxFdPDHLT
yMTWWGYBmXJf35XknFj/AcpQhWZUN3VLaqVwinGcQI3uzsXwfQ+v6+PMzXrSJzo9+HnfXD6oSK/d
4gB4PEORK1cwwJL6LQQEF1HJsOTNFM56OXeqFcR9ItjGODPnjoHq/FBqp3PqphG0XVhFBd+/57aq
D2USOsy29S9R/q2yhjcF8Y27+No+XWfYlgN0n4TwMb0aeBAnbuxgIRiBztL8PvtqdN9c3SYsM0eT
HwjM5EpcnsJdGlWnUJX0dMOyNU47dRvoYMnAfUclzbcCuhCWZJHA5xa+IA+7uas+2ZiY7JH3tg9r
XW4O2OLC+xxyRaPIokkxd7KU2rycDV6kMCWSGi6z1Ss1VLoWNeOKbJY1Fo5inWLYdN/T3e1M01aF
+Sa6m/4JQq0j2bVbYa795vNyPFxm3aMpmzovTU0famnw0q9biYVvtrMqRW7Lb5yurfpYf9aD/Igx
AVzDNcXVoJKc8qLk+b409ZZheBsgf/jtPEdSMB3dcIY3++4aQWDwtxPXPALoV892bhudskXb6iWn
tTknyLBGl149yF2DePqC8SH2wQnnuCYc/i19TVnNARZV7C9rSb47eATzWPkWZ6bPt4ViAQK2z59m
lR3/TgrI/OAf372OL73P+clhIRB1Bhq+MnLFX74P1h85Q3KrSP86+lA6Z96EHgg0X7OO/EdyMCl1
K07mMCB27f1K2Kvvj344rr/qvaJJ6ukxuhSakBAsGo5FJ9pLN0GsKmtshO3zCLgjda75DiAttkGy
NnKvBhEr9em2V5MU9M8tjGyl1F+IcKhFoHilHkLQ3DjOdkgZK7KJT9Djb6TlHUVKk+GugcZBY1B5
qL7yFN2QQqrSmQBQnIzVfVqeMRKvAoIG91tUADYAz7AZXkka1ilY2hzvXGMIu17s3d456a0b1iqr
yo06tLL4BfMLQC5q4Nlk2Q/DDomT3hCe3VWNNZAdXuipDcjEdfllTu8JsB/VLfoqrjljXl1AooUO
eAM9A5bnLTLr63dNWoig7cbyd6cxBAlFC4s9HoTLoKirvqUmgEag8ba5LsrMLsTHrvbtrBK3kFHk
t8CMazAdgvXxECvzGfewIWZ7s6Rd78EQUdy5ykXKv1e9mNRx6OmAAoxxqnYV4aDLFIbjNQGxEEuV
ewfa2ilfRktfDZW5dXhPAI81htshCPs7zFC3++L3X2YC/0o1X/v24NSTsr/rTqx3p2wq9DEu1HL9
FKyf8EJO3ETWenTSevCMUjEU/GSb9PMC+qbwAPnMlV87m4Rt4sOSbW/+3hd8/IE7/rfm1E8fsbo+
6art0/KgyPZy/7kJ4Zs5HELbcMdaf7ITvuzjwwV3GVbRLiF43r7IqVcjhxigPDGFEY6idvWCXeoi
EHjOt/ubO371SIECdSJQ/Jzcmkow/G3jqtjzvYwF6iFUM9gXxTk7HhlMZxZlxGbct5+MCY6+CYYW
bz77owwpIbzbNMqVKdT7b7kiCejvyK8fEQUFZXwHQJpirDZ/6irJv/2lMNnkXVQhzhYTu+I6Uxil
17ZIDdcdcTNJx3r6xiLHVjIc2aRZVdyBnhkp8BG8XyV0QtPcanNHFs4uuBj9nbc/Sm4hEmjlPW8r
P+XdTcLfYNmtaLzQBfdWkvU3hfrH8HZtEE2DlguUZO1NS0XdHS4VpLrf367n9Pske1pXSvQm+b6Z
zUNX+mBEIae0tnWxqOQpUIBYAYi8qbmF1lJneFwue0C4pjRPEd6mJ23+GPM6DGRWPZlCTYdh0gPM
hTrWappUIh5TdY5SZLau0PYafCQywlMX2rLRaK1Db5SlDf6mX2+LdaQuWCb+e4HgCOIiUyc42sle
Ct4l2u9t4Os2Vh9pLjk1wyzi5bU+L3DSlh/UszbSxX7ybGgfZSrxf01YH+NAz3cygsf0O1rc9qfr
FEtmuy0f63E7kvd9EnScSQkasdFr/WW5nSBkHCFTCExYZwtxv93rGgukV8H/ZY6/JooVJ4Uh6fZ2
+T/iW2ZGHZ2Uo5VTFQsbftugU3R3UwUTYxoLFGcbwWEFbnU73MP7I78guC9xkzfw8WLl6Kw4YyVc
e0/22WCGKjujelmdIs0Vgf4sI3jY682hZpH3wDG5a5xZdDR2p0L76j6SvLhlLUdm4zL5EvUkf7/d
YYTqrr55KKK9x6nxRKnRIirg0SUebhmj8ATVMTY7OhMzq6CYugFGOafH3xCTWe6mz1BdndzGOhow
mpz9T6jBhU6FUoBp730OUY63vniN0TXeeqVGP1nEUXHOkfnklmMjlGpNhh3w03EKZ66aDL4iiYDq
xH5+nb/DdpmRmlRNAtcKB+sTl8epnMYP9DmLGYdskhZDGDNsIzpphaqQFkjaX2ohvX6g0UuU/2Sp
0H4239uj/cy2QMk1epLuldDolnKQG+FqCXF+d8GB2tIrfvynC+z9Je7mO54rgt14BM2r8HL8z+Nc
wxpIyldycV/5xhQIA6sbb16h6oAyPeCbZmXXkJuT4A60jva6taeqIOGANbc4ZmdCcLStCg7kCq7I
9rtX6pFqk5Do0pdjly5KDy38fnVoXngKejZlIlPWml1tg+1n7i0hOBi4OqjShCmFbExVj5tag5y1
UP8KUIQ83IUSM41XE01xz5JDb83Domr6qYJzE1Cxuj+ZkoujtGklhZXmb/x4tZQtoasFNbohmAb5
6/WG1xwTyhgRTG5KjPgkmwbDoOL/MKyoyM+C8gUzxRkWQMzk16rXhAl4gILxomJ30m/8a6D/PdFS
40Wh5DEs+jXx9RokLt6VFQZQjTp/GifgR3bG7vqY6ARMAeJZcOLaaLd9XNPHpWULr59h8g9SUcxA
byzldYWSaBe3lJvr2dn+MzofrYRde5u5gUW2JGr+fQm+efWxlc02KRHvcy0HD7qRVg1GZ5+tZLiT
gPevzKz8jPTQKiLRshTM0R6ClovOQKDDbLX28LUEXztoXlUVFfX1ctGQBf0KMC1+VpI9ITw4OqVa
ATg2MfwvqJivvMiJRosGv76blGoLyacT7s+GVkidzU2FoczNyTVnGI6NXuL1elIJRGMKL/3uurU4
f1fzCuIGCcp2AmG60RIxqr5tOmS11/ZtZhgW/a6PcSejUq6f3lObFwu1PN5M76K5pbMzdcr7po5B
ROUC1GMZeZ5ncADnsM0HXACyVqFmW8jBVqh4Sn3VoVPdSMEoxveYmZm1PDcFC4Llt06lWEK2xv5k
FiH1K+Eww2dIDPD40Vena1OgICF7t5KfIY6MSiWG/gf/+0yNs+wwygPdYTIy6QZWeW3NJt8tEy+F
llqijAN4pUPlNzqqjqEJ4iphKLObiAmDv26t32weFoHbPMYrbio7df9zETuhAVKUS5SpsKUwMHK0
Ug6iems/JRxaBwM5vFfWnJj6xI4YOemlRJbFosG2N4NJPCHaw53xbVoRf9loFIiWTxR2JfR8blua
vuFf2Z4jXcJrw02D9NL0sV+TR+DuFX9OaSkNgdPQsnlOOLSHQiQrmhtQ2ZpHXoJ87y9uIDYaK2l5
6ZKwffaw3bq2tjUslfJ1jc4MN4A0LEv4JrKiR38+xTwold4ZksHZFODMh2vkNd9Um5kB1vj3NKMS
sz5BMX5CnNVNurZg7nFbseJpuQLv3m6uL2K6FLtgQi/xH/zSZ1O/r4hMhY795QKXFPAYTOs8MY3B
KlOQxX2F2Xu+8+NoxGoM0eGwVfKw/+zfszA9UkhCSGsk790+vZ7kMubGVP811cwqMPgRs0vACIlO
r+3NYhWrgtPLv2KFW5IPxzcitENmM+rPtIF/Z5ds3ekuTXb1TTZ+qzBhyvaCGhWdzk14JN5ws5p2
o386VPS4LLlk8n31yGoUHvBKf7RYWVmZlFM6DZBt3UO9G1uV4hkun/S4ADkDxR3TsayXun++DLSR
UVGYOUkKEzR5a6+zQuETdrgM3DLmvAoMlqnYUAlF8BufSnFEchPZVdiD19PvQBg9QLeVbdHypuOK
lQZWYYdpwuEvUafyt4C8gm/04xmVnWqSQSruKUBqtmzS2ECIRlK19RJkXV29b7/yx86MUo5+r+Wt
8CrooPozBzNiwl/UtZwbk2Cz+CBG3KVpdXcMLM9d/Mm2wWQ/mFfbqqMDIZ+zIBi97kT1xb7k1Asj
Pdid+k3VM1lutOwaQcYZXzKX2gRyamrvZ+ffb7fxRX1tc0rPMBK04pLAtNRLRRHmOoDdbyt8sUD6
bxyvKBFJTEQVM0FkzNgUXfngZEMWrI4PdUMR1bj6qTQ9ptfE3L2ZHWxsGPHORIm/jJ56z0A/XqS0
K4UUcFZYVYPGm9rBJB5zFhe0IzBnc2qrYcQWqGp46Y2OJXeeUYCfD3srVa17vFNVapIklLe0yD5P
7ificm1Nr1tHVBHUo+qrjT3lTLW1afo2G404eScyIiIqRHI7BW+cNcwHVM2vZPzo0TkSA7F4jni2
h2JmbwKb4i56+hJALRS6kpqRfjZeJnlUeXQe5ZEeEFedzAjpyMUWXiwZ0SLbvsAE4/17ECJpxJOJ
OdHimhBKP4Erk3B/vX7tlkO0Mf68qYl1V/uVD5nTDUC2Of7mVKJBKU1G8GCqO6KqME4RFliIRn4p
CO0osccxS/OP0Bw0/b8pwNpoOIBfPw8gT7vgcgsR2phmeltw/lrpp55WQgdgszyaB1oHhRny11Vh
lnE8/rZD2zxluj9FIs673BVkPPjG+DEs0sIcN6IQ+m1RPjpcsOLJ4LvUkzShp26jTso6JqsbVRhh
WamfIujAzPn6o8NWrW8uSs65pL7KYT1g/BxL1ykqF+fFgyIDCD/xcHQTU7hpGl/YuErrG91454Am
KKwFB3zfBTdyT92iWF5alZ78Tn/JroxSLibje7ABwpupy1ytuTdQCq23gCQMtkWxcDI/lmD6Sn6F
Bmeh1teZ4wZlnlOYLKwhcPXPf0YaS/R22PkNu/h6YC+an6enbFip2dFWjz0bj/olWzRqsVbbxJ5D
aZjRmRudldlQYgAImS6u7xxwRcva9SYk0kNhznyKQtsjlyKdspYPoG/WTwM1cnzgMeUMGmLUyw3p
ID8TLQ/0usc029AuFMAQLS5xKD+zXrT9xm6y/7fsKEcMD//gaZt9IYrgbLHzhKDMGRzuphwgzN13
eMYhANnLci6PpWjVMBYc2M1JPCKbrqaiqOY5jCWxeMeHt/vwg634nln6KTiS4wZiR6o9+ZUOAy+5
4ir8ObMOwKHIUd7XVbfLjGNGJG6fitl+pa3oEF7zh5TfJ73otSdPac2HPJA8FduJazwDWLHWmOF+
FUrFnCkJXybDOBv5n0/mPVMa3uZ9UEO0zgu5/FA4zWKR0QbmX/VMypjajy8h1TOWWdoZGpQuZlXB
jSSm8E/BM8TeQrl6kPCjY11A+cm2qj3Sk/n2dFWVff5I4Ax0PlyIqsK95pYmCJTCJHkwkJRL0tdt
y9DsMHDj+MjM+F8PSPiGpH46EsZ3r0/6hECyadGCpV0EUVw/In1xniS7HZo/h+8XhBdcRQAld1NV
sVX7Hu7Uzrkrp/qvPCdK8E7YkN0AWkwrCGKDvIDTRLObHnvv4tp+Ry7V/0WcAUag3tQexoU+fFVb
HLNR5Ip/Oev50h95j+fPnVdpf5gFdmS1QFOjKAolAwWgTJAqvrhrqwUvb4rbeMVqK9e/FuZ6nHwW
1HsGBxJSkU+pB3bLYp19an58Y+plAvY6m7xmR6iljnjonn/j4d2wiUXZOHYXy6d+DjwuOkoXI+CF
aspxW+eom31vH5VgAKUKbpC3wvMtdTGqyNjhrB0gIR3t0qGnpBSf8nxLFhSKgwPZ2yI/2rGt16yZ
m4jzABXbh9wyzDD9tjb2ILBsLryT2tV8eB/ljTq7Ka009Q3FWWRiGseg7hbIAmlIMAU1gyLx5dss
igDzmFtMc7S9DRE9lbsRp87FbqSvnrIhuxRmQcRvpa/1P4M7fT0FDUW0IvMlal/zw2Jk9Jbt9mk2
XL086fqUm5eRwB1GO49O3b/yw5Yk8e4m3YrJr/spVhTUnp7gvv8ZIRLMGp1l1OSrtlPp46NocaP5
HrAHSYho6XHsSx/o3vpZi5rpYwTSH8l51Ai3Kb/SYGSuJYuDv30CaWV0SuGfcMiPt8MAncDsCRzd
jpGMOsuMgPVILRd2fzZQ91QHbjwdH59pxAQvW6aGM+iWLqlpXM4iqFLojPStJTdyu0zCTjf0265Q
1hF6knQe9tIiYHo0jOE9TMHU/StIkL8/2/FFdkqOXdsmy9bfFTpPFrw83zbQyPcabiitClpk8RyV
SQSbO5qHtcOF9273Akcis5K/dZFVOiVZ9mmWzDSmIDmrYxBehtXIl2KA96md1xWgPtrrwTG8DLZL
pW9uwZKWudSzKNVpjW30UBEHv08ZgkowtwbMJqAFoQo7UCqPQLLhcqC695kTVzdSBkm9kvAl28Bq
hjyFKKoUxMJLwe8XMX1pUT/O09XF4GDQwS0fyaukxPHvk1RYTXVMMSgq/GtTQdvK/Kgw6O2h/ydr
X4o5SVjcN5B0V0jTk48j5AD1IH/x08C/qd0ls3cYU7YHtZPOVJnp0wH0ObH3+zWfjQF9zdA+f65P
kqUmi6bWcoIAAghAVRMvtGhV43FCKekbmYbgu9BDSSQY5m0rrCURwYdT5TUa9TgoNPU0Ugn49zln
T7/jS8hVYOb6BS7sNsrwgFfNACzH4nvSGPi48Jhc6w89PXTSMPmFlXSqetG2UtZ6TXVHGlFhNQrB
+GF8LykgqqNf6tH8fiwKUtIFMH/cLDPZqHemhOk6lRKzwwTrj9NNKGt1GnheDnBZrydTges9pcUi
xUQ6Y3yDiz15s0vbIIRsJPFDxVKm9XZIhVgjq4mouFW9Kuan5FJ0r80uoeEjSkbBNdo/Jd2IX4a/
SuvX7q5Qm6Z23Cxc+bNasa7GeTkv7lT1q6JakAQVaNrrKSnZ0XTQzsx97+ZlDecYDXcq0o1b+c8A
omoifEtihuKqWQKNEo8vF1USxh5M3toqAv4vuUqpGkYXFbwxOvvZLpKyZ6auHmjWRloOmP9oN8kj
R1EYHqMqUZz7eDpRC44khkzs3505YNqbrxymRT6YiGocYIl1jtq7UQYhGakPyvXt74qdRJsAubbm
0NBkpDafyH89KoJlK3MQlIpERHshfrQtm+1sNZG4cKOHPCvveSqIxfxH0YDpZgVYitkAfYVH6s0Z
o2Pzcl8veIsqSoUof6N36caJCL0VPW/dz+EoHy464gxsxlMN71fN62JaTV8jLRBukUdT+z9Z4Suh
lpy92cEBGKRiY+lE27vypqO4JZ0r+x6n3CmeAs//BGV9rIDstxudyEgoershAvH9kQtMGl4Jd2oB
TCmMoNKvJxxsd72QZkOb3LNacVRMjtyw2FB/qVIuPeFhsEHhAyJN5UEKfRUzwK3PYpUgOXoK/ke3
EPzU6MDB+uq6cJ2Upj+YPkXv9oaO50sB7em/GI+zE8CebTR2YuKpnHfmg6nS4Mkx5EUMeYZGwVNH
sJN6D39cYxxL7L5lRYtzOLo5KJgObZUFQrcz79FYcbyVADer2OfPmDQpdyKO3stdVgVygC7jqvKh
jjC6j5Vm3mQjpGf97062ajBt5yEhQ/5TB5M5YG6P3HmYtXt304d73Act61iTdC2W5xGQ7QrVpZC3
iCt+kkt9llVgb3A4g3/TUK7//V+nneji5qzEEsL9+vk70UcRn1zd564cYNUeexbUwrwzlp1Y6QQr
2VueWmqPXCYxg575G0grKCrmHnqSeqbdeOUOPQOJjDDJIKhqPKvbZVRv5IaYVRu6V8lxpHl00Za1
uXQj+wVbAVIdka9XbBWCAP88mYq1mCqFPc8CFjJISM4eEoOSlcq7HN7LxgjSPvX2K8/sbZfCvvhz
Gx6//hhv3aYkE2K8ZIxS2PpblBj/9r3cX8STkbMPql/DTDAv7Q5LI8XhE5rcJZZtxURF8HR5Nc6j
/orh0SMgJ/U45cvALGgetQcGmPpCjpYrfDL9jrSbGdtZW6hkTgfoul/F43IQXAFqrauN4wHXxczl
pLEiAVQ1hw73AkRlScdeeSjxvcttZhADxv4ciVVDv2PyGZxd72tWWwWDTUN7pcYn90tNi03efDxo
u33jptT3fhlmZbd4xpIGR7vZiYkC+rRQcBQ+bIkPVuw3yIMlQ3a+xOkIsjat2qbX1A0O2GOKuTtM
4L4IYhipeiElUOw6YrvOZy1UrGRP6K1dMTtMMYKOi0EK2H3Mc36War2t6kpfiHjmWxC6bPaamTrl
xc1XI/mHOP/vDe0LPKJK0ysUj/dLqf28bMCDe6md6fKtxNDZcDuI4c2d0l4QJLA0dKFrix8vxJ6H
3kL03YblvZjAk7+1LM7EXlAZ/MBCHhMXHk2M3epAC4KYCiqHu+Uu03j0flsIC3iPXieYCHuWjFet
z2AtI1IthGll3InparFOOszNpXF0480TIewlClFESY50bxKg7u6LbaG2QhRKM5Xmq1vRc1VhnCZO
r7Y8sSOicqWla8XahNPhSsscx4iI2qH7c4PVmHNE1z91mXvOILL+YoKo+ZUmnppMAwzInMqk2ow1
Mj1X+oYZv+2jIfAnEg2VpX92BoX8uodLtbKqJRPJYntmS22CVfnXeR8z3Gd+ux542FuTYsA+nMaQ
S00j56jY4KGZdMDF/AG5UVipLk8IrRwMIzWlvd0HP2sMLYL0eDL8o6zUg7MXH9vShb3ctIR74o7E
99IvQ9DdR+J+ueXpxfdkngMPMozToTFu0NvjySpoYzo+W9yO136M1zew0V0euPaoLrytDSVZXykq
Y4Ev0gJfYBGllClw6ys5xOVMhJrlVVyAuDE2RofrzEkHKU+XaqSKgTEqs3HmMXE6x8julhFAeR7P
hWzS47IskfNMJI/FsqoMRZAOi1RSSi9xQfAkjdQIexJoPVsN1PPdpaFqWqMXZt+o6SXUPiIOQQl+
Pj2BWX2OPsVEfDZqkM34jQWwbR8LcqV52HSS/COkbTNFRL/bG/FO3rLCoMGjR1U0R0VehTob9bcR
S1EcH2xzdpkcEMO8WmrH2kFG6g6On485ByzURC/0Dl9m7fFpfBApQLCmNL/Ovsby4uInTrTERoc6
sRZd5bznDKHTkdasKGQHIaE4Jomm2NWWud9qnR6FUgt/C2EDVh5tCAYLAjwkcE4loLK/RHVQI8zb
2QgEJOJ+gXxiMTMQkJ9e0ZLdNFSIZb0n5VPQMZJIXDQVZt8rVdTHfN0o9Sw7CcD5kRGW1IGUelyX
udhW7zTthOH/KAwwfI4XPlGl27II2jx9sQlxNUxErhD6lje+sHMKi9O8u+sBDMjb8dh896uohSC7
E/jIPlfTIXbPY1lVw6noIhuMXjJKkCzl5Awa7DdARXC2+21Oyl6srpsiVt1XGtB7bICSTSSNoAdj
/YlWVbsQkLqb2mm1Q8aahCfleMmsr/vLlpN8+xcVfIBrgnQRzsUJKX5NNlGb6+YFVO4G3Oif8oGP
qJ4Kr9MwpBYdv7SDjZfOv7nzf9hnq5GvgM3SobsMQ9l3YpzPf5h8XHmvOM1EXog9DFMlYUPT6GSh
A6Hn4lem1S0durhdYa2ZbSuSTlAVrleliEI+4CJ/hzB6fhj80/Hszici9UsgJEPrKhtk5mCdeFtO
9KIlggTParOwNlNubnM6n07LshOZ59o3pU83T9OGSwyW45euNUJ/mHpVFV1LSsjWlgo6PGTpK8D8
j+gQWFK+ccT9/mrE/aaRemMYEUPM4rwvu0JR+cUUBDJh3Yx/2DJLXKH2k9gBNG8lQH/D4LBDcNFu
MeYNNqoiZfB75aBZekUhA/OQDnLUpXllelxDM1lNzjAXdj+tT34FdSeoRs5STZPVOzlbgEbtQNOe
FJpWJ7S/u2plQ9fsa35TQFz9OrZd4fZUp7YiIUgj1aFCMLwzyL6b1WoqYoJE3WDUHsOObqEPIQhS
SkKYPnQS4aqfv4Ut3nIYFrWHWm8vpGP92k4kicbiUra1Q6GgeJrTL+IFyfXZiC4B6XO4U7BpxUFS
Fb9FLJ0FnkpHzLo3uCbJx9QgPUtnFYPC2Az7nbUS2+YfZnxwdjJlsxTNDGA0PlRgNs3YGbQp+8ZP
+LOQVbxufRZfqS4C5aa3Re7BntfBGuVqaqc1zVsg2LfpacJV11DYeuaOlf5weBTH60gwhLEe+nD0
91yCkxdjAw+8zgf21h0wfjfWm+6uUMzy1EJ5N7H8QFN4dMHw0aoMBuqSwIzuFGi1eVn/7lWpTJrt
flLY/O/C0aECLmoTOBOqy4yPrlxFoB7m7hJt/JfJkO240XRp3SKdcxoN72Uqjp+vLX777EbNJQ0y
B3GE7P3ISAc0YmmTBR9BIw4s4x0vVtiVvuv7ktV0AP6aH5gW3wvmAZPNTnFCimLlnEa1KPkyXnyG
qMZALJonLiG7RexyJcDJ/PvZW9lhPVJdUSRJTp8LuKkYz5vkt/KpUNqiQBpFqc5FFek4R3OYdl2L
o8By5EEtscgUndLFFXSoX9Rf24+rx5opr/QncvowVTs5U9seouzCyrQomJgDW7bXwKvMkqTbDIVU
fjsad6zFxCRG3tj4JuUULyd8+/XXsLeMZ2D39lJH8dJfjie+eVxP73wgzRakT0J3vAP06eesszak
vuYj+8jwRO5P0BP1iTUrdFn8A2lElNuGsgNxP3/n0LFZfp0XmYL/v60K8w+Q4Nf6YCbDlLJmcpM1
nUKQuzQfInAn7fKL6WB0lFeQTu42B1rFsG/77DPOIHy0VEIlp54YwFIqLM2MXguttDTtSfyNb12H
MmktcMQblvTVEQ807oEGgJJN9Lg6QbiCZplnB912tiR3x8ILWlEJEaRAB7pd+FrfEwZbQcZlb+hT
FRDP2xSM1Q5jj153C2GRRM62sfUpHp0lDcYmC5sz2aVZhAYgeFv9AcDM+pknxqg7WpDbpkZDi4pL
tRau5H1zHs3SwMk+W/eodomelcMX6C8Q+qbWS0aM//6CsCxHfLUKaBRfEX1D7fuM3Vdje1RuiEMo
j3SQKZ9Gy8mUv61Ofnh2OW7dFgvFMQc6jmFHLBjV+c2/bpuwvl9dno9/ojjBO3yQD8nrUtcLvMVc
0ydDwOkHHzMKwR6Eygbp90nOn2hnLU1WXnEvQBNoDgz71Qyvs4mk0CRbbfBbIDCGUs1PQ8fjsFf6
BsZTwP5R5/UeKvpOsLgDvc214pHYY1mPi0FsrNmTH+KVr4yYIlUZzT14QiUlL+hl6OisUZwq3SX7
M5sPC+KZeRyYsu5iqnbqSeDp8kWXbDzQ0Px3rUNNLpkrSe2qwYFcgT2E3JpXGLVU2x7kQRTRlBvd
3LfVI52sR2QnrXBlamvBDVZZ7MGIcjQxWdbxrnDpbII5RtNM0+y502fHDaRMzO3DZnQ+ocMeL8c6
L3tEkXHqlQK6OXjBepCKdUHDF6CiNLQTCe4KAEuwQKYqwNvQKchei01BzDkjywjJONmvP/D6Rk2U
T3vpMu7TrFm9MOIPQIrFwt5muEIW6HYmBtM440Gd8dPlWiX/MWEf3rKjoCTdbjnMn8AqlWuGDy3P
gJTNmczcg9Ve95ajuiAKY2UGzLjSjdvpyiafQ/0Yev6hoF7k3SXBnco6QYv4ohnm0n4qkgntq3UZ
rU+32rnfn0F4/qymWpr8UbSC46YsMjhacqN/IMdHUXQknka8A1JU6CERyb1ziQVQi4VWBSCval+k
3E4qI1/PEAUx60rLoGapnQJmYA7QHYP58S+OdW14bKKYAKNc9bFE6dOE3lOqjxKSByetkDw1teXj
osSjY4lVpss+V0vmMJWmznrqf6HiSICR7Ng3UCpZA0/KCWqdwGH7HgXsfBhgQ4hJihaRk9UNBEaU
Iydx4l9Tjqv04vM3I7HVxIYxjeccqbbRI1evJLGZqmgw3KV6zkzvTZzh5owLbUbm/RoEO7JWYndz
9Byjof/dhaUuXNkA2utltxgsl13kDZ5YLPNrOXinxtLafS2R0aG00XpzvjiXcxexUIilWA8Aci40
qYd4PCTcstKZCrL4xx0nV6DSIn6X5MNncdNMumKF2e7lidScnZE8EATZCFrrNmvJWb1D2fhjYY7N
PM51Qi8KE5rXQT/19JOaxnvL7lF3ARkh09l8chfpzQGlWWYZtm2r74PrMIJQJG9p51p+Dj/2wwR1
RfsaEqAr+zABCOuaGEG45DOHR6oKqUWneaI0Kz4grEbgzDqLt9yW/DRIfdLyrnrVPOeHsk3MOcWG
TZ2BKhfntgSVyVoImENk9fMwlSc1Fh+To1JnP9I68hSzO6r0sEZBz1dmMkdYcQ9jUTco7qpkGd/f
WcCBTnKui6KAkR6GYVCbCyEGibKqeM4VH0AZH3N3yOSdwGzeS2pIK+TqimvY/M93MdRbimeD6G1K
nqX9ImdH/taTiabgDOMPn3fsQxxLAM/47QffhKbzkimvzoZCIG54wyyMywb5BCz0KDzjAVDBW9RW
tyn/dETOz+QGym7oDNptjY41KgXw08biRqOk4VSLB6lsbItBVZWau6KOJLVBh8J5QM7wwmC26vEk
eMUd6O7jOd8CAxjIilFzIrvu5u2XDV6GUsGhPwiCOD4HS0wlxvwqeYDM/hyDdN3nvkQVisLsT/NT
vc8AN19jfLfuAs3IKK4ovVHdY+u1rip9UzMSI6dC2fCSdBy4VX+F3K7ZKkhEFgAIZOg9nPIYA4DO
62uscoZqVoOIYS6hNX4L0UAO7uvxh138qIEPLPfV0lxJ4Z/JZ8cn4Epuvm84c9YSeuuHMITh5X3V
Iuc+DB0lEULD0AA7EVk/Y+KJtsmRo/nXhUXa33+VgO5KHb6hD2lteVkrLO1VAsOCyH0OzfAHjMCp
z5GcSGicbWQhjtQ5lFnxuk4zwp8LfFxSyy/bF1dmdmJFWtE5VpiME/LNk0ofY9kwZe0ywB1iZCkF
7rPDq/cYgBsgVR8oGeL8zCT3saWZYRQ5kH7lLlDjhO/iJ2w+MB7LYTVQB7FovzEo+Vc2qzYdaMpp
xmIneUEfmOjxzZM6W292ww950FDoQCpp1t2WEYEzMqnZtTo4rk0KaxIv4hpdROb/yXhCXx994oXg
8OjLEbRvLwxBSBhLS1WE0wleKNJDM/2ejtzuGlKhHHHOVrS4fYElTpugv6oyZYA28ihRpGFaQK5x
ZUmvW2qWiftzZQ56vp/PNKBVRy5ilrQCXpGPaDI13O5rjrTCLe9QrY6FazaMb9i4uH9COilGssq0
60yqBPY3h8OxApr+kZLc6ZxZy7XBB3eaVWKnjT+m5KICGA/zJ7SmEoc+PMlPYtP6WePJ4fpaGy5a
lVzupY181nez0U0c9yZj7sVprCG+h7axJ8EooJodDYHRfLDNxxRo5DOI5GcxQ9gFhZAtZLzKiyI8
a4xbrhn9z6uG5vEUmzcivmhNrUHMSPx0CgpFh/Bd/UqGspLrOMp+T0g7rbjt0D5Lk157IjHDitTF
cU1+BBGvd/Rb33vsvPoyOoVGJJqdGr5d8VrbEqFnUbbT1R3C60TQ7A4+Edw7JLxaCunHph+aGZk9
5Sp3OPsIYqRI8rYIIByhzWJNORIbJlsrv6lSD7QpV3wbOi1RedNa0a4XXvLFcoVP9uIS1QP+Dfi1
FCjf+m9j729kP6c9mVtUb2XaHAoLJ4iLuUq3CUewOCC8QofXE1N5leNy1SOPv1H/vZxdKBIxb25w
ez82M6T/E+mU4fhjHGa+H7NfIEhWEm1Xq1WqA7KkEFEViYZcfHI7di0U1D/oR8HHZjeM+yxMl+v+
Nj7swGid2VXP+A9P2uHnJ3Mrk/I8jyiyZsRhQZSPMBh+rshT6ZB1vfm1tDudD2sDeDHX6V3gIgvh
2WnKK333BXA11N6T1cWuXpXmzolp0csj4S+i8UwmNwYMkYjP7Q9PPYcSI4ZTGp5CuqWl9QTq1xxx
+jBr4Txz7EXnoDh/7hlxfgdZ8z12ITvpO81OQjn+PtNV8FPN9CzXbs1pyCaSvwg3HdB5kRqsiHuo
18Sz0x0qENr42z9YOXKShc1cLNBkuhqxlcqHqHQuxNg3qMEwzfvRTGO7sjEU6SdldmYJ34VA8NaR
blNuD96cwzePfZypEkIZTv3MRTRxe9nj/+tiBPoVLBFQBoJnB1jwPhn3h7JpmLfbUszxDWdO0XCB
9cRt0R0ddiUj31Y716VhI0NdNbjyLImAPBpTFTv0rImwYgZ6hubzfalJSitiAtBOItzmM4huuGAX
FMipGLawUeMhi0XeMpJEMvjNEHG1Aeqx1578Jjc1f/tReLFmdUoAuULs2rSM1QJEe/gYoQ+DnY2I
AvyW6z2nH/4MiIijX+mwP2QBmokIuLezwY46YKx2dtFjyhLjx+rE9LvAoWg3kHj6cg7GkQb70+oI
pdr+6wkwG3qBhV6smj3Q4t85W3giI9gETMTAs2gtFtv7qw9kXXqNYU1o9umHjoshI4+XH/Ss7NIb
i1/ELXIfUdtQPXpzoMqcsWexjJnZp3B+GdUPZf9j1akNfqkcKV/sjVD39RY9i9YZ/faRxVRSbUwj
UZL68tliB23mCxt+E3eY8IB9lN9eE1e0j35JHDVIN4rbYdcoFxzN1vjD4lY5XyHgtb9gLAFC+F7Q
EWpsg7/vHAzLYGlaua83/xeA/TXHKrKp7Yk1Ym0hw3nVyZtIRA4RUM1Hq3Rn3NlqFNyLMlwwZJ5B
Ma8TfnGn0Fzb17TdSQA/Uh2qwd1UBonHcIkCeNfc4UaG8tdOLomHn6ZQqvO0oIUi+q+NEsi2jubk
7vDMQV1mcveemI3iu4a5DttH1z76Mad28HKZ/QwiFBNJzdf/pxDAbqEaixv2o6plZXLBi/wKvWqg
SCVLRglSt950pUHUdEOv8e4EaMzNgb8TJxcP4GusMzZGhNtxMugo7AO+Abgq3eOAJT2uYvcj0I7V
G4Umx9WlHd19MXSiEtRerHOAkTP9bWLcOgf3m3BllYhmQ4IeLLMl153gDOxd5dwlHfk2X5KKZjTj
a6lg2ulYJRN1wZ/ujuuW9baJNfpIOu8h7tCnjduE6qYtPTkj40O0odD32W+gJYEKU4gZ6PjvvNOo
PZOFprxZusqCj+H7iFbF1gJ4Qt0n3EsbqB4bppy5TNv8ciO3Dl2akWBdCYwWvNGiOnxEZ4Szr4xk
vwn1TtYFCGa6oo2Bc5ZiGGJZClGaRU0CrHqJpb27KRePwvcAj2Gg21mFdCrI4azHN9UPJc2qX8Ie
S71dSj6j/v8AD9KPUOSaVI8i5ImKX4Yi8AHAdo0QGDP2JVIVM5rgqfpv6uIrB3O2/6bVkaN5OG14
npffE1MUjxok6Qj+ETEY/knPfk1xJJl3qJkDcHr+A0sZJOY+aUrQVuE/bfZoimErDxzhfyUmsk8q
Myt1Hv93D+i6pbL257gf76dd514k6ITWoVUIXlHfWOW4ALsT8cqO+uk0/EKLWHsVwTa6zn52/fG7
DBmJKEzlPBH2o/Xbs0PrOSYN8KDUrzmCvKUwzA5Kgv/lmKXUk51P037yUiArpGpVzoou3x1bR5CU
B13qlc02nBPP0YLZ0+4I/nk+roqym95KJ4xdM38saVRKeQ3i5Z2WaYrE7OCBX/TFMts85YtFF2Sk
xEJAntP1xXi5qzxNt5cj0yw1cAZLxtEyMczLsr9+schRvfqUqTghZ1lSr9/ZWU9/TAkfbuDYgkpa
ft0UZt2TeOI85em4Ifm5/4BqrmZNBJqpMXb0+NONfTAx474i6hksgJOoIdL5D6OyQAJP8xl19zvr
jAC5eJoGid4FIT0OIAWFZy5Ufh51xfjSwhqfpTG9f1jPZ/5/ARZ39AeAwSfSRMqMSaRqXrApxoC2
aZxlkwt7Faf2K//iNo7e6ypLsgJEQielevwh2DQzfS0W8ixI7lW083YM0eChJrI0JVG9FpbEFJ/f
jRuRWUdCITznTfCxY6TB6oDSEH8U2IZbsH+W4itoiOgw4Rlj8n1a7LKnC1WsIALDgx3HtuhbCmnZ
W/42tALkJcVG6l/Kj43eIvo4dt9/7ZtKFxx6uEUpEIMsNzAW1hwUjy4It1VO3/TbV1Iit0Qkdf4o
ndUsjjQlAXYzba3XJmPIs9A95pcXazXbY9cRKoGErsCiRypo9O5sYdKBQmBy54PRpN/U6ch8oviE
pJGPtf3Vc+sEtBSYZxwAzhaOdWcLd8EgYAoGz5i/XROBTPK3Xvt4mNGv6RnjPYyO/DyAq4C4GimG
ca8YzQcNiwxvnOKwSLaB67JpTOkrgR3X2ipObBosHoywLveDVJmbDEzgsVkMWS13MRbnkuWcbWvc
fYZs7WA7/NWKCVWCFLyiDbt+NOFa4IKQ0lIPUe/m2hNfFIWyZ2mX7edoewuK3fSglbrFHRsR3XK2
IgFvwg/q0jhIrggyL+hmtdQ6qoHt3IzfkXGmgquKBHuKWDmHbIigMPBJA6CmiSo47OcMFd/jKFts
9ul7Mh5td5n9xFqVZdHPmdPIc5HDwOPJNDhTcWmlfliERSNzbF5aG7ZPkbw1Y0epDJrDF89jBgbB
+HzOd7ZVv9GDEuRoi0GTSXhOn1y8Hf2GZesZU+JvDJ/Er1tNUA+zexhqptypQtGQO57CqMVPGVpj
DTt5Fe3HtVUXQFhuDvnZ7IWMLpZrzGX8Wnc2jwNFDWPxOl5S1QsN58D6F7ZKRxwwZHS8Fy9COO+7
r5Dzm/ioXLT2uzzTAzl97cpOHrllE66dUctV+P+O6ZdVhJpUT828B4MFzgGsjuIUgHjPYRxEuvlp
1vWIE8r1hW9byDf3/OMw4spoKLwETBvtyzCUnW8VUDGTphB4kT1DRPLb608EkC1HxLQyMhiSxFqV
vMemSe1RQPNaXq8lNf9EttRTf/bK7VP2rYdtlWg2W0Nk8KLBTAzNrhlCVhaGmVCtr5ytlbApRR+p
OX04ATfYF+vRa2+xUxRC9dMp2LLFTiqb7U2r/v/T2RdUC71KeeYLF0dWyzu4TTzp2w+MZBgZ+m17
+zmAdogWfslhWHedP2+jo3Ep569nVpkdRDINrwASvam71zj3y9jJPFR0uvQxpyKU0lPuS+sCCKan
sXrmvHPbW4lRqca3iWi33Jwiu5HeiLVGFnUWxPC4vyFJWiy+RILpQVGBCe/ieau7WogBEnPfdLKj
QvoVfZQXx+jitNIaN3J+WDV+x/rier5scMigDbbyz7QyXzlFtwp+pdUIXfc/UbPM02LJ8WBdtg/Y
PS2Pnn3pUb2Q2KdQu7r1u3bAfbe8r9j8z+T1fR8XI3D8zKEOYKhKATc9sejNp+7QOfx0unvGd55S
LBi/7JMUzMbWIZqU97ixt574eFyA7FYuW2Yxflw41rClJoX/ageHX7bn2ESpLwZGDoafMVeA/VFD
Iab1m3Yw5BSCXH/xhi4sJN5jt8XVEkSBwqfQ4rGbTOMNzP90a/AaPuLW4yq/MLru7FFjzgySZFTh
EpcNLObh63Lx0np5ES9uc6F3B00Gh/a76I0P4Ll/lE6kv2Lz6+0+PPC7DQCyYSWf563MoEMiftWO
M/YEWM7L5wmWu6/fPa/gptGDpTVhuidJLikPUnHieuqj701whh38GW1mhjfeJ5efUxL17LoiCY93
1CiuA5PK7FJLCYvmixiolw1G2GuzsVTxnvFE/bTnpBvV74FY7Qc9VWOHaiUEQ92oH8knNXzjpy8v
RG6ri0dOGUhIsOewLSMlagq9Ml1EDc+Fw2DmnwiVhTykr6K/TCAa290OqoHdJfbYlKEzcBFftuc7
lVMi2pxT8DU4ReThPQqCfAHrXbeIvOXDx/tx5FE0N4w3B7M65imd0Fd8ZINNVNTPZlu0F6TR/U6D
yZvXA/NXXPBUsoCHbgQUqbZCh6tZ/aOFNrwt7Q1ZX7QEPg02gXa1CJu4BjnzsK+UJpxQvniEkzez
zVgpx1gfUhQnpRlfWFf2G7G+5OG7HJJIRmAbYcszlxKKWtCNKYgvhP2NOxAjvh/x3+8N/sS7+QZy
p2kt2EhsoaGn+MRNZPGdt1W5Orag/741+wBMNlQd51ZrLR2Ib0HXYIImzqNDSpq4N+MgZlvu1ZN2
q4L5aSNXcap9mYjy6N4CEclXIMA2x872lrvHwxne02cYUmJnTeUhfuy3TBR2DiUN8Fy7HHEN0KM2
HQyMS7IxKrwxPj4RF2c5pqEWXU99/fpn+UZeypDCNiRNt0pKVg4EEHZrl84jegV2nXZXqsTrcwFT
VfDYV5/f0FVGmLNRKx35hoabxmfuqsvhCFw+3tIds7doJJjsKiyKBdqXZPNcfkJAeZvcNmPRfMZH
ynGHvuhmFgIKClffeJ5lPvuvoujS11W3pvO61Uw/+/OZYJN4Naw8qDv8yGxasGUBSOCwCcd7Z4PU
c7B+9T2OxRxjeMKzZhOonag4Da1f874xFNA866BOOL07+fmdpyEBqaHTbdl36P9WTon12bF9dSkk
M9fAWKH6iRDShAtJErBnCAB9ylnMWCBovEm2c336vBoVKGEL/CVlm6zGP23NPgMs7dvLIRb1e7yY
50LRpj5yV6Ln+TSrELA4puWRUClFG8M0qIKEC37fRtMzVNCcwBbLw0hK1FDaWLDCiiufo46LulwZ
4G2K1GAMPz3U5GbCYKvEXgUjTOKnUJIZ8zXz9Pi7RZlojn4yBp+225g4qmzdC3K9mnEUgAdTwP5e
eksKagv8A4plEBwRlCsuU3pq/Qetz5jxOu2Mjtcz4XBEgLeGzd/mX/BulI7+TpGld6b1hOQWnEKJ
FXjJWPDGcejSA6H0xz7UVuxXxQSuin2yjxBovSlDPFVCdjsxySc3xBwufx1GtfsfI/g7izdHEbPL
Q4KiFk8SqeMRShp2EfWUHk2nxaEc2gmeo9OK5MLxZBvqR9XEFw+GjnCb6NSzSwQ/nzHzcpzurpUu
MrpDMbnf4s79pRfqjNCS3J/ZlZDNJyGYW+MtRX64CkUBC+wvJOfJ71t6kzbGeElz7KwoRajpW6st
eMujXNuAE20MzrUZ/CBxGzP5vK83OexXtjEF1BCwV+5l5RqATRX20yHzuu7ESB+B8uduMaOy2BSD
nVn3F+koc+rJIZLMr0nNM2pyk7/RKSZe03X4OYwzzEtQojAz372vtwLqkZqJCijXhoLrq0cyO6af
d+JRKFJkJJDn+W/391Q399wMF7crxfTgO5w5JsXOqqEqqBMXHbSrdsGOT7Pepuv4jFtr3v2hi+hW
k46RTEiB9EdOnRFhPRvVQu8/H7PYdYpBydRw/g1EArqJEbVhW+hLdNHciLnRNcoFP15LksG71fSv
JxQ3Ag8a9PB2esK0+KTEIiEBJzw8AFitfL5JN3lIJ91xvn4vs2F4yFrSazu6KmlBdssqZ/vhWRJG
pVfma4aq0Asf0uYWnGd3DAODLZpO3s0vl0oW4sJcg9+N09+pCq7pPv0NskSNnPEOv4OoPakyE2Xn
5nrfqT9QtL4uZ4l5XN1bevveye7+fBq6dDoGID/zrH3QSx4WN87upDfA2GlyiEyYlyos3OA1qT1H
sPTuPQKx1CmDTHHyDFnh2Z4BNzeLJ6IOHZqlvAxxmGhDoE38AI6xU/dtb82OfuM9WjJysMwGWnI1
/ElwCh4NtsZvlX26oKfPH1QBZboZSv/M1UmpxUCSjVxZFVD2WWkyjT5h2jr1Tt/i9ZBUFwhFeQrY
vuLSNqqjvqqhcZi+KTSLrbpTLZtUfPaaqs7lsdNqkFW+VbXs9GxXF1mKTsRD04tB1ZQvbubCb4eA
BjdQATgnZnUcH3KwjhpkEbKkSj8bcznngIjzZGA8RpRoAbqU+Eg+vQdgdqQpxsR3JKe0HQ4enKLQ
nAhHKv93j79bBdpwS2thk0BgXo+Gw0gKSE8gRh1+HBQzsRalPup3BiKJN+fteunXxHyJOVjR0joZ
ZzEIIqAQ5QkzcJkqxD7B0UXEpjaP1LxmK+hnXA/hiq9luBzBVg3Bvgni885LkJ4jVNyvK8V91n3D
oM6b2u/jASVw/IDr4pukBroR0EjsUPa6T8A9nxWTyOcFFBxccQf1AWwpM+Ewnajwk11WHUqd+AOn
Dzm7d3m8oMPoD5XZ2Er+kd6GOIORW0plQ+NMdpimvMOPIdse9ARqC+ASfcJnnkmbI2dUbe7wqRot
xxhU3SZXjIBfpOUGoaR66RHiNtekd+17Y02zunPEJJrn0rQa047HSIqx7VziES/FsqeACLFn1XGz
Zwn17tIzab00MY7cB3CkKCdotoksKBojwOcov5Pt45xn7wUI2cReNgqtrkAhzRjBpIpITdHelm7U
w1RIXSKEZV+NB/mIrMCJ5Bv3q9YE1Z49hMo6ayXd2rc4bzyl5Mo3fkPOmbDwRY7dRQbVz2ThcDS9
GUgNKuaPwS2//g712dXEDfD5T3ZIjovoWIV9LA6JpRfAZdSRt3vw2vSWQLDeZXjZXKqbje17fUpz
m0t/OaStpnEkLyf/hzg0a3flIlz37jjvtxNMaSEBSgwi+Uj2cEAYck3t98QQjzoV00XSIDXVmcKO
ElQEy74YP1qyH7+fW/BPk4LtUz2lbuwe4kEMkoE9/jd4ZE968PqozBbGx2FXdRE3ktzxdmnB5nTx
mPO213muJEE73+WzeISOeHIzcncfUAsgNcSpZVkzA9wo7PJ+7SzVYvAYEkW+flmZ5R9jiFJ/t+vb
RGtIq4RFTy/Bu3BwSQAO02JDuIrDifbxVA7O3jcJvp9/JcN49sW+5zAHIXyKawcefNcw3s7HMd1P
CwMB1FrmAEIhHV0jzJT1HBVM+nF3wOIVWa1LrbGdyihQr0dt+0q804IXsJ6iyRS15Vs7PndVYexo
tklZwnexl198npknfBnQLb6gA/p59ppXQAQCmq6P5La38Llo5wTt/DGU3Yf9GetrCFyTcgBNYKHs
jisW+5xpet57DtRTfNLAJul8Vgt37fmDprck/iI1KvUIj/ZPvzLb9beGTmcLwm1tdup8418OVWF3
peT4Bk4iTrCVXtMg4XbFmolPMsbHlDrCn7Bt+XEbZFYH7TbyvFgQAKLv5uWWIMevsiF7FsVokUyj
8UdjfcpKidA5dKSO9QhzGGekeJ5ybDyiDlNqqMriMhCic7HMcmoVgc9FI1y3JE4T78otM+OqYfZs
+M4MasL6rKwb63i4Aleg2DM2Kt7+9xXlWuyp59xiEmJlv/PPL+ssbaxHT1aYDjK0TK7at1FbWh7d
wa148YJpFn/Nj69l/me0j4jR4fq2AeNsKyFn1YZQt7KQOklTBWHyxO+hngL2wLJQsSe4zst29rdK
4wPAQd1j3XTHWVsHQEg0ZDIn8E6Fr2+6W+y1Otp8cQlZVgNiNNEgfCBN950rWoS1sEZKwqCBWUyM
hThUr7An71++XZU78/UP9L4QHAcRdFeGw6xC9Ns2nFOkkNN3vZv9mtCbUiRIEE4eTLRlKmaQIkrM
7LX2ZUbfX/XzqFJOZrFeWfTULrrbqWtj0GoTypl5JEUjaxJj8Jl7KDJaZiO+yRGkbuQHU9CUQvSs
MVcVwCBL0Y0pmZotMeXwwYcT6FxoUZWwAsauYwJNY7x1DSQJMSO0LTrjGLVZzBwgGrD8EofZJitJ
2QFq05a+BxAdzUGAv7I/DFNzfarzlD2k8VCx1RLsJoxFjxZaLbtTJllp4Yt0fCrOIv29IbrL+TnB
a+ZV+Of3qYp+/1zHWFVWAn6hm5kBI/GgI3kyCxoFdScg5oiAbKuxIBGgP3yov9QMoQWX67UuDhkh
PsYUrFWQaISvLHo0TMEZ3+e7glbHf/c4I35yam10yVDlNhXADulPpF1C/eGskOa8r99u+SE1ouo4
MpaFv+qTYqP7WReZVpPOXNNg8EpxlCayyNs0UcJwum1H1SaK7dXkxSH+fed92Il/WBQs+Zo9Ibs6
AM+QB1Nz4+1mzAxic0brkYDLyqaLjBuyUwAh37seyMy1O/NddFlUEzMVgBkXpT01YqnEpvt5RmOS
Ql/u8DyDwdqPspLJeAdQt/VjTTk0CrM3CUj/1BkCfVon7hoWkJv4GTK8uhIBnARZIqLFjnSUkBzZ
temNR7IVbvJ28h/6TdeCOrrlrsr+zeDkzzVis5Ev5Os7EH58/6nYcGq090rpRZQzF/cOtDQHzkmA
lmwWu/k/1jM2yaH+i+xtYX9CizdYSp1ErwRDQh1Yi8D8QzHIC/uvYisVCiS66PgkVKbzZTcEb8pQ
YNtL04vqMrEZ/F7qMorNF4He4x3p33fIlSL1o551NHx+Zb7plDbfe3H12NpyB5/3goxkbLu4nvc8
6S1V5tL2FYJ3WXpaiPmoBVkWngGQwrOjF/nOvgVe7klB0no0IoJnOKpErzQUX0ER8sLA4DNATVBV
70GFnQ/VnfuxDFsiMid+3xZJxS5ztLdkoucENlNx/zF67HfqFMprgmYGpH1ip42ifJG6aRjNhBS0
PnB/ZQQdSSJyhjeCd+WiGC2pw0C4AbJJUnu2EmGD/B+k55QOjcToW/4SwlQd6FkXVhI8DBtwFcqg
NN0PSxN1i5fF8rj66mDYxxcfDeBJEJ9qMRq/dYrSqJ8Vx/MUzYb0SyIAaPa7uAh9FMJ9u0Arx/Rk
rlSYUXakfN1uYX0dlnbE2CX6MD6Oz/CdlGFYtGgHezha9vcBtGnCgka8NWvLD1FyEGRoNmqck7E9
SmiS1iScvQkj3dQ6SQhQGg1XRsz1+NM4y5KTe+Fh6EVMlMOiCK7fxsFXXXMhPrHRniTNb+XROJVS
GBcuM7PdX5m11oYbk+SLezq0ITp9Xcu4BvA099T2PpY08gAtcTrCtiW2pEMCzk3uaO1qeDwJBIqd
SKvTDlnpsQ9HcZjZqvTh9oXCtkJcTY3SHFSOSncMNAA1tdXGMGGFJkSRquG4t15Rc2Q9G+La/ptl
sh+s7MwiTO1/igGH9UE3pn3akybkX2qcV+WK2wavXjobzzsOdJIQLrxMPVdxrEDfgTOiaKbVgPxK
fKFwPHZ/XSpJHUacBQFXpgKiVdw5leGjRY63+WJZGtULftGbUp+ttTimoQ0mdy4+Du58PWOyw4ha
g4hdP0sJNKioF5LQ/H6qHMHTdugNrLBbPPvKm8ZmbzmEXGICI/fg8ub1fEwgO+TUCzbkyhV0/GQ7
HZlG7dkFyymK36nXzZsc5OfqqssS7rWe84ReyDQNw4fO2+xK8hPoAN9B0LjJNkPEM/uo4f8kMbkg
Zx3kGvCs7pSgSu6NxNfWK6uuo2LOrY3wFWvNwZJnQNFXndxvraumB/M7aiG2MjIRRe4x3GDtZmmL
EGmF7kCuBww7yIHP/FKfuF9IqrjRZeFdKM1ktnjHHbGcv1Cp1/kX6e3ihjfLjHAWdzmYdwyTlZnh
QBfDU5h4+OYaRtq6FOo650dKxhM9WBXtEdtxBXDemyC861aCjX5v8G5MTB4V8h03PLlNTMpCZFPW
8zGe2f5Rw9XJ5oJYDq3cS6MHjOTUjzKPtMb3OHepFqlpegtyaYgXjl2NsuVPQrLlSivwUjjxPcHm
Kf6XvgjMOhfNNcDyqEckwYreh+nZ8pHHiWbbw/k9d/UNB3MSDW9cliKptmn6VjnhHXX/G2heUdsa
lR4Dwlr3OZ2m+4FbAIdhMzPtMmmX00f+qmOLXveKl++r32MwqHDeZeHgr8gkQ0dreN83rJ5bSpA7
WDMRE50OF7fkua3kKLDetqRohAN1novoQE1Xc4aLTEiU4WtXG26nkyKl99mVouzGZC3n+uuVvdmH
CqQI7iMAJc940KtzXU9tqpZKguRiruTHupHvLpCvdpg4awUJ4AaVracqK6YHP+rAAMzAQjPtaIQy
UorsCgP34Eq9pl2ydTqAArMxiAn4nliEghk+70qegarkE1JCUjMYDxLEgizoGjLvZai4lytLwG2w
jcu6NCIj5jfWnTqasYTRVpzmO6zZ34clhqRUeDubHBjR/Qm4COc8fftVy8/7v6EqCvbyri4qmB4z
NuwqdYpuL5XUgci1PNUb0ZhihLBYDnUbhiA9lBSCScZjgAXUJE893bVzLDV+CrL+znDXc4koM7uw
fgH/gSL/uYP+NB27GCnUGxfg+7BtPjrThHF1RPJa2HAcHpZ8veNvLY4liv1DmfXaYbtRPiI5eHAR
1GO2IbfR3OzbtK1CPpIjimw/P4J6T1SN7bqAZT85fsTKa6QudNaUXQbHezTNGg/ATqzw0G3QcZSD
bKbh1ao8AH44sEDScO/QA+2mfrX5IYsHvSsnKkGETHe2b8VBoFiPC/nWFyG/7NWIP+OVy23xuAiS
L/WPj/xhg9iMOH3/O06PnRmsq2xS4intI+3G0U95H6jSud1B3dEPmLGU49pG2OlynB1tncwi28O1
ZqTFCR8mQ6NLTTaebVzaOrblOAYXZGUVqB4A/E1q3nP5NuKJrfb9x9LMUj6VmMUniwLlsGA9q29l
XMs6z13TLFYztD05LsCiGtZlt3XmvK3LCNhF//LNq6c3zdkOLXhrNhgncdx9Q0lO+G8yVLTe+YrG
5Cm26I1ieffk9lpaC8GcHckqcHBdzJ8yuglSHSE7paPa8ceX5VnLwMrQq0Fkx5kXJVKvdVdwYeXI
YuBd0e7G6xcCJ0FsOhOI6170sgtK5zU3RnR3QYy3y0eeKCwKzGN4CnULz432XsUPCdGOwU9ftBeK
yi2zS8/3iWnzRFVsZgIfedUHLxmeBkJVvEAdBh8JWjvIePXEIlu6YT+wEUvRI3rEzDOmzA+++alb
tUC3UtZwKPqSi0E/nCWQwgt+jCuq561frNw++sq+PBeeJPDi8IuGIVb4nWaUt4/SNROwOtc9QENr
wzwx97XMUzcO1YstKcWAQquQSfinSwjfRrfBIlNkUMMW+FiNU0cx6LXbLfMYjNKeyAI1hCif/8Oe
uSq1knRpd85PfdFO0/WDpUJ0pxdSBtMsrqIkJk4kngYj3NZZulfnO4yI1zYj7xgVNlZk7zWpkdIW
2quCYc3CcrPvW9NGD/0j+7Fft7ItKuQbxNreiVWm6KiA1YQVG3BW3dpXG3lQOR1HGqSlWDSpAxOL
0h3HNu/HZtvKUhRGtCvvtE30pnD9/V425W8x24ID/8XbVWoabohG2haiyN+IsqGGuXptOfNjSsd6
QwYAd6o+ESSFLXQiVnL4W/665dog5XmuPrLwqq3c/nJk16S16MRZ0nPIvauL4KQQw3PQp6Bpi7xn
hVLWA/JEdRiLf+d9vVfWP1hf1YcAccjUtex9ioeJaQRYAyPXnd+0TPwIiPpW0LzAG4PBHK+arhSI
fplGTQQLqUy3QBGYnbNDXiDvVfxm6n9JSOb4CITjaqjoCLM3F+0673FR56L5r/Eh0dGDtSELzyG0
z2r8skLlWm9KkdQbqEwMQ4rQG2YctxKj4wo9LxKCJq7Iu1N+Kq2ORke0SvXhAcnC/ji9CrReE18s
4ME0rOp0VHJlvqkjrxgop/4pf6oADvEN8nimjYrPDdeXvLmVWdvdy+WYjLSfmFNC5hi3ECkTRob4
dGvGibJNwb6HEWdaH6WsaCpgZZLkI8hk/7ZgebWNO2wDlqNoFKblOQOvrZJEmCvgWNMxG9s6lujT
onfHqPhW9SodokCL/fhW4IafHCXRA382TxtSPDS482NobhKtjtGYMEsqrRnfHR90WvSExUTBbXJD
FWTZO4hfvptuUS2Upe0G/Oc7oBKid2KMZ2hAmrfwE0qlyJW5bSyBEDmWd3u8/dtkXozMl6X8OmWK
V4n9FZ87nTrJiLmwq/rzSOVypKkxz4vXCAwaD4XEF0yg5od9BivkZnp4AosEutrE3zJ3Lq2uCHwy
BMp++3dm/s6jhaaVBJZddooPJXiva1HAUU77bBLGRnkuuiKIhPLV5suiPRU6sp60+MRVayuC14qz
jj5lqU7u8I+6CYHsTY0e20d3hVfcPErJ6JpEVdcOWzFypKh1o9lZf9Yw9a1bVTiybgXxkxJs07m/
W0S7RfyvdjfQe9576kMGs56nZQah0ziJB/4nnhSSilMb/xp8pCFwG3GLgJQthejubvVk6qvBxu5D
GoVwxZ5lPVfUwZGdkwZQ0SCiNRFK7O8fLxp8zLDdtkr2dtU/8PhcuZtpGmj3Kh86+BEE7/YeQUEX
txMUwLKr9BGjj62/dXFp87xgoiqCURe6zpWiEIeMzu+gWrPon4B0t2Huv2uySSWJNCbFA9f5xbkN
uPvWLz0SHrwNX2zwaFOeh3ctHlRps/YmKzijvOLkhnfAixkCD2Spz8f3gKaiVZM0GrdzKDpPG+EB
bQoFvbAEuEUfy4CF4lUSOkX73Y5EzcTCh0YqdaKt0mKSMWEmOL3W9vpeVRg9bqP8Udf2JVoPj5fg
3fAzcw63dCWwSNMteqtKMND/JzP3KdYuhUWeMU3ELyQb79vQorqsZypN/PhayVG5LStFyMCMfw/G
J6OQbmGZ1nKNccRlWfrwfVxRPJkoGIKzBalGTucMxcqV03UV1KSuyqucY1NNB/PcTynVPRryZzgo
F3L2G1t1J+NOW25QzCZpT8k34qofeZNuZkv8k1weDKgRXblFnuTs/Mls+ykblRyfGYsYAS30WAMB
JtT0ise0k5fBpMTlSl9+kGdC0wXfL0biB9rX9kMfOAIe3ylBD6VZFGi0bHWbXh0qOtrlK/EDNIJf
oSHFeA1TzSc1RY/TLmG9Y0De9TPtfKFdUSabcTSTzwteBli7uKpQbulexg5uwEbDMhNNjKrDU8Ra
/IZ/6YIW/iwZ03c8Td1x63hos1WXvMF4t9YxK7PYQrge80ODfbUBnFhXS6bnIxwEFt8s7ikWCuhW
091u3tU6GO5V0WBWOVo1pHimG7KL2HLtI33fC3zs56F0WlKRoGkWqwZr57fEwQ2rk++9chs/O+CI
PoNRbR6CeSKwyRaQjGXA4rB/vXyX0/qb6Bbz014pfBhc4vDlnTGvhdc5E/5aelARGawOtAz6XUbs
I6pF5b2dDu7lVY5wkTX5pH3DyuGmZe8nS9HLlgsizNK1BeZGMLaYO/Yip5hqekCkDn4R4GcR37/6
bm+PDQ64x/FzVSM2v5/cu1obh9Vywjdrn/1zuIKcikRIx2R888PRM1bbuZiDvj5QBbXL8SNrepI/
cIY7H4DXKyYUEkRbtKlQh+KY8meX9bNKIG/ifKKM9oe7Y5eQXWdwj3TDIk6d4GPIjb6f6iI43XA/
BHehYzFRR2Eo1xoUQEtXedFe67OOnWuU9V2LcWWRVhAQKhVBatrxuWT0aXq/fYnmBTby//bBOPbU
hBdfcdiJOGBfFZtYv0SQg5Vw0XO5RAq4FGR9JFDmFUMq5MMjt7/A02fzZ8Lp0c9zGkceydJJZJIm
fePmqVHbFUXfCnL5T3i7A5XoY+o0Vh6hqjvkQLi/qzNKhFHsNMJOr6va0njOyw1pfQatyRPc4vRk
cWFIOY+RKYt1Y2V3/9EfkUJ8q5bjDEFBJFoFVFWUpJ/inmhzHkSkiO5Qy3AtFeObIHGXcXb5tgQh
DBWigpypcH/DutCk7unSoMy4KYFPRBTENuNdKHbEQNlid1TqIgkY4KBogf/JPjhM71AbE5vuDJAy
T2NEcZvp2+Y49R9HuFe64Xzt0EEBgWfOcI+wrtXwllhbLPgp1E9P1m0btCbUQ1tOwDUpFOeOh3BX
I305GJx99knXXD8ofMMYY3cM+clXTbBwHrftPPHE9qdu/4e/BKuGomDHj2eEaB2zXGKac/K+GMmH
LpjUlGjYqHhGUUO4SjRiNtjYM3orBLzmedbtu3JUHaUbv9GAXIWk0FZhAk//W1AFqLXQRhHQ6Ibb
Wc2GAozh+FpfMAUUhIkxELkf8E/kH7e2ZveS2lHKtssGhYGpF1oYNYOzekZ1B2cjzQkFS23ygafw
QlcMYuCyL1Zgdhp5JHY827DwTk5xSvW7xbS+bqTWe+Ck/lq4VSU0xwIT0XHTGdf23GZdmymr08ID
oznUzomYnkQU9Puto8O3OcW79rDpT+Iz9hURYmPQV5XGtDjuz7PSySf7LdhpWsiVgyQ781ia7I4m
3QyqdylPYnL6ZwNMEjaqjEwkQSiCOMHllsVCW3sCCx83YinY2h+WxUAHICZAOYQqzBfIXhYvAEZ2
nm/y0No83RVm0S9f0alTGdPaSJknk2MdxvO3MgNJrZmZDGkriDH/agYiN5r1v3tohYYnYLpdjT8K
9pjyo40PfgilPL2qqv68ARdkKaCukj1kVWEYV9HXuYEWutifz6vA+mXcowN9W2Nm2N2jCjBvChFi
SvFQu0JYkMl8s8t7mrlSRd2YOiqaskiwl7yKiqScQzwCA0mkwM5ob+T7ifzvb8ALgZi0qcGsNZHr
IsBQksXmJVR2wut1VoaptAxgkkLAUFrUT8VjOkpG2Wl+Vaq7/9fX3yAV1aaSmasQHrjA+IYRZIrF
SD5dnX+24h59TryEcB8i4RSCDPdpJiMx5DDGVLUptUrHfjUcEwDX4j/BNKDnGcGyZnOYn8PTJdde
FZnGvd9QavKEztSoGrINyK4eSqqtttqgXhz+kN7po2FW7nAswdWiD9f9XwbTJ4LB4vuoKXELtOz+
afhemziHqBjY87qCTYbCDM+O+BljHUvZdyNSgB2WRj/4Vd417+OB6jlVT/iesqBm4DRJ0uUtS618
vv5Hn8ED5gLSsUO8IHLlHp4DQdJgllc2Keam8oAVrLnk+3cAdqlnpIuCmbz/jFUm7MpcWDSTHDT3
32MqA+Yw5NzYtVaMX/KMG1Jq/wiXGhEO5fYMT2Ol+t/xyOssq1TEDfALnKTa+QQIo7lZjlZj3bTw
dH5gdAoLF34b02JYDukwD8fJx8i62YZ101lDr0AgP3iYA/E+g8HXCQR743lvhqA5ZDIeJZf4F4tP
IG3VfuvC3v1X1tQu7MWiXLwCjVLhkv2BVVUHAHpjNmveqcJaO/lRXYJsM8btUdSUAjv5popC80Wc
l3D53q6E/DfjDwZ9TjQCKYPfxwvTJFlEtpHu9BwVbF2ds9+s/9OJNGY6o2G3XqP0Vxxty+IRSG8J
a3aCkHfuBvVMVp1KU6/9i5wGNab6kL+Y89kU6bxVKv4i490D7zPWPLbVb25QCFpBkm7+i1ZUyyLX
Kkwle0T676zrjEjwiW0Qu7MGT9tgLCEYh2Xccsj5gsvJQwQn0aDnVEzqPLJAxwJbgOrJBwXZehUc
n11JvMvzsgn1yFKerizpHKh/B/7tz5mu5GKJvZSBlpzU2mzbSYZ1SYC+9oDKW2LA+sAoVaRiGRmq
BY6K060XRMWu6bPMDkSzce8CAFktCUFmS3yThGFye1Ejk0nKQ5QKyJgBFeTeSl/KtbU1yYgGu0q5
auJZxdYnF/LoCcxBstutGJ1Ibmwx3J+WkmCWWi6t9hA26Ok3atchymEp1HW3QvWUlxlhzRawr1+n
H43ORy1Sya64aZUYzwtVE9c0nt9ZjImZkA5VkBTsslHQGUSdSgYuKwS4jbt8P7AJSyO0qWmZ5Ol9
zpbuVZyrBeJw+P4aRtaVOgXea4V0CtVs6M2kX4XukKgThwXlcJdAJ3SA6zttySw23EMNT+h5uQ/2
xVoCsqZfD708Lv4IPOAfe0OXprWqr3tnvk6eMcxXPvE5n7dbzB7yXZvQGtT98iVF8S2HOHdDIUCN
oA+fUQ4mNylIydRpJklFmJEooCNDWXW9M9CFT3OxbRYznBKpmzeyvYP1wTkKqN13kLS+zSPdRZnL
UPbyBoIK9BVvHDULeiJQ4pwY7TWCQgKaOvK3Eu6j5JZBTTNnIuoEyYiTpAuNLVYoR26ucgkgPrO8
KQOfJ5DHbPI9iHprHkku0hdyXooigh5vxVJXSKbKmLd5CNSH5uQtUVaPm/ss8XvUUWYj8xr4+NYP
siO+EuGcykfvNZmkeSZ5AVm9IsgIQ76Ux2XRr0mEZX6pdCttO2+pqHy3AxoK0vVIIX129BNkXDG4
7LDChf6ZzeKYlblSRlvD+sTBFQkwih8mhb6MryjBWFwxjO306VT0Rq4RZTkpCBxE1Ud0Y1EPBx3B
rQes6a4I4UU7fxGEDZWM08GMc0G9QpNmp3A4exSExqeUg6QOJvLkBAIUCVPtg28jkPzdeoNXcOQa
2Z3nm+OYGZGiyvzEcwI6lBY1eN0hLLm3hXWEM8KrqXDKFRseQnXRCPazV4kvXSH7C3nUz0jvl+lr
rxijZriRgZN0w+AHl4wpMEtePbFfdjRr7x/MXfsm+r3J2we9IXWFYd0cxjgMiRGyFW4utYl/m7bH
nJGar1LgwCXCWlGJTgB97AMaNnqkfN+aCTKB8ttKkJe9NGLjx7c0ax4Iytd8tcgd7Ip4My4mgMoA
ULeEOiUCu7mk+uZ/GIU2/s3KMv+ZXJryLfqZOjMGEt7L1PMcZUQS0frq3+LKpH1lTZl3obsymTZP
B+q6NeYkJAQ6w97NQjbSPj9lLZhPST1CX9/UiVCZ0Jokt8HiMP5OX4jug2uwMn6btupLT5CWrB5P
ujcxf+4tkk7cVEKZAcqC7LiZL/4moDD0aYrZpYWbV9xpoLudTJ05KojUE/Bfi2q1E2kBpCVRDtls
CDg9BjHlYxmwr0SUYwae8R9TzJhi0mELrZCmhPsXEvjWo8AT/ExKa2dV32zh/7DNKY/kFTyUjNQ1
HIHTtgj7Y1vHXI6Yaz116mvHBOTi1xyRicLhQYtop37afbezLVcfyQ+Y+ZpOYXtW1Z3wSQNihDUT
f8BZwo3h9dRftmOP82xjWS8ujWLKtQMGnD5cXjFU7uNX+a6M1P9IY1hlLy+swDNHP/kTQt1+gxsh
b5PehenLXZdXBwe5YSUbjPxEwbavv7fThWeAqwa2p/epjD0554xGs3JbqjcgJbpSEv1Fn5QCsHUT
ZTA6aU/U1/Ma6pV+h9rrE2QQD0MzFJ4Pz3IVWSQkJZJzZYRRXnykvNWva1KsLrQ+LayIQ80b0lR9
4caCanfLi3D+RrOlFTlxhJbZNmPP/Q9ljsrO8LJ9yeuS1lLYj+oXfr99ZKIBv4G1bFG0DuFhAzc6
6TJviwJ5oet6Usbl64vhmW/CQ+Q+hrDTqecF1sYqVAhbF6sP63/BkMqAKeaw/J9NqfKh2W81eM6J
A65fjtGfpUaSWr+kAbfddPeoRUBRvh+mCtvoUkScolJqJ/HLQppwrm9rkSRch2oWUtqtaZALY7RJ
S1My2eYFa85sGqqXkqoNqnHWVDuUrDSQydxofc4jkeJn7Sn9hP45NWG8pOnsQ5XlhuRuSuWgAKfh
dDQPUQh0lSkEl6y/Gl6cGdQgDC1CzNx50Y0WiUij30xMsKexuTiEh+9nUAzjQrwDEl5KhQj/cBmA
xhPnjEs4qMp1UnM1dKpwgUHqqi8f9He6znb3/CUY1iBhxGAmX2nEy7Yid5iG8A4g1qETfyqdIfVb
SxOyOzzkzKryGfqMg9GqF94mHmcTvMZ9tuXRwuBrW8b3BGyreK5OXNBqormxYB3DDmU7YYnBpdzc
yE+y0P6jjbzqQt4sMdqwDNGCECDNoKh8axrRL3Pd7v/9iuCSOB1d1Dfp+Ap4m3HEqdH3x65EkVCl
MYzRh2rP2C0/CrT/xLwGvM+ZbjoRPHQ7CekZWF36ccZB8lpQUBLNnWp8xkicQmJtej9xkXy7PEID
XhM5dxdTz1IqRG1QkN9QTGmqFBHQvoxaTBQPzSqZfggC10RHGL47OQcJ2O0wgK+FkTnoIj62V271
kOQjPGpX/WZUM7DDgoWHJACxqGB5Di03JC8ikpIwdICeeCy0U0d79sZ1a1XnEFuvzW48oEf55n89
0oJbepan6bxjAmPcjCXwHytOiBI/+4t5JMDkpXYjAX14U35hu+kA+f+gEVuqRObmf4JJq6jyoqV7
F70Gvgq+ie64wNDOFqSexiyUSP8/6UvhIjyVcdDUDRZGm3ze8ykM1YhWvHeqIk/XDr3qhREQFzqi
7KK3GNw6Mp1dofEZR3+NF9/WEwg9ic8WHOsg4Oamk03HPdTAwuNk9C9Q8BTp8Jf6ClJlJz18I9Kd
szMlwQC41/YEueCfnO4nvT5pJiTPEiFsqElZGrFcir9bVETc8z2tJBOeI6y6lI2G+QKmT6tdtrz5
pGokq13WqsDioGUXKp72dCWeEqOazYLfWBvf0QTwpvIWuOl7eWexlfMoaH8HwfohCHJ/m3tm9Aqg
aJnGca1LJ0Lk4Bnew9dZO0O0BP+DEgjvGHvjgmSeoHbUMCtvR4gQsKHNy72tVs49OD4GPsorAQe4
xJWTECVGNXGAFf1Hrqyl6jlhml+Z+twWpgBlZWO29OCnS+HB0qTLsmOEOC8+zMrJkuDZHRuQ4UJk
9HHfR22BQNM/a+dH35nKr/0bGW+jHft31zrosAjoFLuk5PqO0fRsjN+FxSAlnc04rx5fhkHkBjqY
uUnbwz9HoascR7lNv/4gBOR1hIahHr3Pixkw/VdzbhfNpoBJ6dCA5LLRPN+vYFr5tjsWW59eaAFW
jO0wIglR6a3PtbnwAabJuff7DetmsiY8CMAW9ZUf6TA1VF8YWAifaLs16VhaD/3Aft2DZIDog3fp
6pSU0vCsOrNrUv4p2VXPc7PVCJVEjOElf/tJcmvRo/qv5yETGobrtDHS7dI3xvPB0MjLSg/re5wT
JKjU5/MBfBowD9Xy3jHdTKODDBPXlBVpepvPWSvBSAKo323fT8qLezk8xNcjgXEGW3Ru7VuJN5Yn
U9REz9W2UBphZ6rzLiNh/yijC1eMbAxw9n4sjzijbj14kj8UrrjpnRB1f+CGzq0QnIHkWM5tBSKw
q+QzbBaPBb4AUtUGCfiK+ynaPt/i/bdK+X2DYU1ug9DVSIePRZKxbl/poydJnjeSn4/DUuaKKq2J
EcHalyggW6m68mhIEuph35m1FNp5y7uucyt89huviXQNjsFiR1RvykrIeX/btn+uFcfpksZW+uEW
bPOqupgm5jJJ5Fgq0keuvh9GFTHZIFrw1sf0zAyPe97Rhr02l6X2Eif+7HmySW6TgTCTE82diq+9
NfRnYe0nPrSfB0ty/arH1JrCrUx+AL92KTzjqtkva+zT1BGA2u9uUH1MSNFan1uiBKyXPvTvsBRO
q1ZsYmgPpjPRKJKuhSQVOX29hAdT1U/sz2bZAh9418bmuN+vnv/LaGM2E4x9qxxzejHMwx4ukqqq
w1ML8O5fIOvgK7mQYyv/nlgY/iKf4XWxXhUrj2MjNNmo4TqpvnWClID8LVccN4TmWhqUloRq0QCO
ZjY5hXRC2f8zrO+zERwh7rhmMXLsrncXuir2l0GZ+UWvs4qQXnAo2AJT6WGogXqAAlLFUZA88hNb
0WA+7SKhIavmskRIlclYyPMGULJdxjsuzslaPkFbWWBVZLJiapMaph45E3XfNSdOYLnuN4QkLHsI
nvce9+muZzXj+X81dJF8IlMi9pYLG5ymUGC4lcQr21yH6qRyAX0aUlI8qe2/OBIynMe4LU6sMxP7
dh3N+1e2OhFZiO9xl2YgKBSVhWEo5mhK58qqGQHiVw3rGI8ZY3/t1PHY+R/4fKdiamx1MCQ03Nmc
F4er7g4qPVVhXxf4hFUMeGA6oLec2XyW9Mcz9y5E2Phq+3bSojBPVz2WL+XA0vGDm5h6ybsprZiq
3TDH3sgyh95jvFyis+2+emHs6eIacC2SHZ2ogT+FV0/cJFEE5skg520AGkLP3OmE0s/srBR2XPhn
qiBLFZ5jDDN76KI8JASVxwLWHZgQlnhzdyTYAtInnOB7pKWNSGM5OAZI51pPPAJztZsaInI8Tvu/
1m+VyjEH1cPRLa0B0F/BxiedGGYfptth2ztwQbyOpgYVqcngTIfNWRVbG8kZ3r8G/JB6CXHcxNrr
cbIN5wL0jBwls54uCX9OKSW0mgtFswRL/FO8nq1LVBpWs2uplNdUUw4ldQVmgIA/dgBkITsBtsjS
LFUQoXuob6ACrEPaoxCzYkpqwG1EcpUZsSMjpGSEyxWBzD4f95pBE3nhJK8rQhFdvwrhdr4Hx3u0
pjeAGG+NX99af3Merg9aYRW+n1K+NzSwexAXt6RBRIscLiJJDQ0sxa6qXaSc8OqZJV/qGrV3EWXp
UK2uAEFnCeZZEfUSFoZkYbz8h6mp/55NPB8MnJSUmtfG0p1HcsIsOD4qSBp1VIFjkcE/I6uMA2SO
WNdTMGKEtqav0hdmYzwadUHvXUWOdg/ZoGaEfY8eD+MUguxa6SWCNn0IMwHAUVNOkS9nc2wT8uh2
bRSeIchCTe7yyCKfORephIMuaMjlrLb7v1WVn+4rxhcPXLMosSUtQH6tULPSNeaoo7wIvCdN90OX
tP5uk+DP556e26Ne2pQFX0jYStHdgcWqru+PZjRj5gS4YyVAh7/4I9RdgzkEJZPl5A7cxlMR8DK7
HfTSkkU++Qm4EkOXimFsP65QzLo44ZJXLzBBrO5rg32gGPZW5lmFLkOmh4xlv4PAJUdlEMR83RyG
B5T421MjJR2EofMZ11WNWavuebv/2gOzzbJxYiutZ3Xf9xyKk2KitMUbvWSnxeZfKJcsmxB9fIxX
AB4SWoOnA0rj5f55CG7thRN3Y7MZrrLJJV1eyA8BQOQ4OhJ05CIwi2agOd3U1wBV2E+oNoxtdVLu
Efb2MxYil2wihSVnfWIW9yEPPE+IMYS0nFSrvuroA6kqcZnGg4KB+DklWLy9p5/IRj95difI2aCu
GqVK/o29B0dAe0HKOzsVEouyDE5C4X6kyp+qa156QkvYjSKsWOYz/bi44xHZza4fa97/41zFjPAi
b0Y1i8LpDzHOkKgkFzmkOmnbsGqHxRoDnArQbLYPhcCllzdAy95vFzl4vojajsbn+593j4bCQEwK
Gr5i20TugoAUhCKMB2PlDjkWw8Xv8XQHEmDc2RS6Bi7s4wfBbsTjwPIX68A8bBkhETArUKxeHWxu
sI/8IKo3wQdfDzuckkCCDOmgS0lllo2wQPbhmG29Sz2Y8rznoaXe58vgfdFvVcewkh8sQ6B3/1CU
jNnmL6bArDtKCZXQFdio/G15f0+ektcSwlRGKBlOAB2B+bgRny3hECtmoUpPfEdmN958z2mK9yB7
fST1Yhp3U5wP28VV10cLAFnId9Eg4lHNelOR1bcrhyHeLMIB4tBFqKIP8fmYHMgogiseCPzFDSv9
6RYHz6QW5j+AFQXQ67NVjxaVFOKTJYRT/NapXb1VWgn1d1lYoXpNqxwEJ46cUKqufqEng7M57Z/T
EBIJiBOu1v5hWzYnPdiY/IFupSZq5QdCurseqqdk5e9E248i6xP6GKKqRuV5bxvD3N28KXQY9uRj
PEFtrSmNgoNBKnz3eNk+m13TOWltUcWMFw/AqB1s0LoSZSlt7l+SZe/UrF0sK7NbqMUR8HBPKX2h
uXb3YiwlzNWA7Lxt0FibTPo6yqieVGKTOSYfgHo4j82GCPhL/6ue0E7B7E2+Svx+SNM8P8LlWVg8
PLnSDH91mxAOpvdJV+9F6mTt2pYJRQgOFpoL2CqdxbDE4qSEgC6EVY4v3Ku+0VIckvao79Y9Us0o
TcelHCWxHxgfZi204SRles0+Yfm84ylsEzDrU/r6GrMllVgq2oCTOnZ7oxa19NtfC4PXanatPGU0
Xk1/YTtpAKk7u+sC+5KcNYIING+GhKIvRXhoVMudPojLLmS5bCvjJfxIhRMcdKFIZuhWc9UA3cA2
KEfJIQIzghPL0mgbjOvBqNga1hm6UhnjivM/leLbL54MDL+i+ymGIQiOavpAser6GgT8wAaMSRi9
2p3Z5BKUmDFX/h6nmGY6sHZsmafPEBsk86/i9ybxH9bUuopU8goJtZGlQnB2JbuOp/DiL8qoHjzY
RuDeA9UA4SBDSOb3Jidt43EtNtXNU9NAniAb4qBn2iTCAgyvmwebGt81AvYKROd4uW5kaVuVzoBM
nVPLrjaOEnk5mBTkWesYsKCAIyiGsuKwp4167bRrvqtcMWV+r9EUmVxINZnggr6sIXUKfl3vCBRd
rUNAIIvGtu2Z4ZL4avBzidBSp3UdOjPJ69v5/lx8VIVeXPujvCiIDyYIyteqcCMUBvIx23IbDoLW
tBg8JGu1KpvTBr3O6Ief7bnID1jec+kyeEavUJ0IgGzc6bKaOJfa3YVVRdYIIx+QXoreOo5jjfYm
qgLIfPraN4FV6AZ8fCxk641uf8aiS26689Y4ndi5yPWB7gOLAn0epbi/egCK0HYvWfgoZbO3T5sx
Enhf8e2WaS7gG7qBd/kKtFOWVI4DX3QfyW6V7jyIHcDNO3rRj9pyzHK1HmBkzxnZLgvDGus+73VX
t6ndvflYLjwBeLV6cGCVvEph+e6HCaELNopf+tEicWGLeQ9kUU23j+M71tNVhHKE6HWaInHney1Q
5dKyyiX0QNu+1XjDvqGhB2qNzrC5xpeh1pAHLn9Y6POnWadez8ZhJuEZoLBJDnLzwM+7JgRIA1es
hLBUt4lYTqALATR/dRlHbKR9iQQwqowwhxS65kK9/wLPP0i1SBMr9MOJX5LIFUuNFkbrDDLdf2kv
0bpW56V2AKaV/v7spwimQxge5aBgm+2q/G5uVTloug2AMC6gpSLUI69bF4hwVnmHeZB6uiVWZ+qx
aYUVkgEM8yOusRsFyEKGcyT3AuKG93VlGSXCDkPNDyS57/ToXiP383vXsaeUBOGYaT47bCgjzg7M
LstUsKJO19VTPgaRencDENb1duNtzcVSoEor9s0oM1PnA0Yt1lhQ3BDKq1acLWmuFDP1AGcnqH+b
X8D7UG7RWQolXG80g8jqViTSNFvum5kVOw7WYjfCegs9/jSSE5LwNRYkileEF4M/5eRzTYAdOQDm
7syESdMiaiwzAYgRZXvrag6XoGbp2jbndRkTAuK33CfukjRn34ktZEOwpxV1YwUf9UOv77umuCsx
wI2f314kCJrlXX/yqs9NHkAY7ONc/BhfhvcB79prYHSRec30D6Do6/nRkEf/QbM5jjI7irKALOS9
99SbJTnyw5Q6mRA7KbBmfRmxZkbh0RvYQ6A+Tlb0Fj6MUOieJjc5MQXMFXIPlPoLJUrv7pm1FeLd
VhuTd95hmb3SNd7ciRVV2nrixy7/sHHvDkV0AtZ57jUqdSU4wDJIBNSE21Q7GNvCwOdX0K/A3biU
wLVFHwMOgKqI14A9gokrNAUZE40rUrC3KSExNQzNn58E7qM2GgDun8MRCD7OByoFIv9Cmg+70R6M
5VVZge2MM3knDqKws0TSQXy2nncy6NkjwR5hzx8TVrnylJ8cR7HRmMXH/PPoL5oyY4txvQe1Lk9P
1gzkSi2AbZXyrnkYjw2nJSdUfnY8VlYVY7XPgDGYuO+zQ2QsIddmWN6GCSrwHYdVARsu830GNfX9
b9TTCio/VEBs0KrDpSr39oDiTlvQ2Yk8d7zprrERbivni5U0MHQuSJJ/H0CoGyFI+3/8Jc152jYQ
CI+ZiokejIc/2a0se5ok6kvEPE2gsEUgEHw4yOzb8eYZYAch2nxFm0s1t2s5K0XSu8lO+C5s9VWm
H1lYDl9oHws2SjlYp66qTzEyAHnRe1eFoyW/ZM/2hA7b3ZQfU1QE0e1S3paKPDktOxhwILKJ26tK
YHIB+TY3i/gyiYUi398eDP+y0l4Pv0/x0OONfCY5N5x+57foD/gzqMcO2dh4FWdnCO+kQS18LyQJ
hLE8IbYn3V01Pkt9b8dm5uTtUXhIvS3BZhJAq1CJwWCdrn/+1WvJbvFgBmCVSJ1rZvJ4fb4cI+aR
AnHpDUGFgB2M8cZKLdCoGpFtNlHC/biczrPqEqk6pYyCNjefPCiYwfIt3gysXA0Zcbh7JcKN3N+R
3F710wpITgia8WMjN/bUEt14Z+q3xe29wCaaNmzggAZVmyw9GHgMzQKlHRE7DrLLtRnSBMif28RF
75BN0nJY7/N3wP4F+Yqr+/yAelqVbfmRoSosw6EcFPc7wryVYEIggIf2/geR9YLtqQVzZCnqtyAt
V85oDD3rTqdUNov4vi6CougRqEZMGCCu5IqWhc8fZXdf8sQIKr1/41tVrK4z8re9VlkPThBqktAb
uIiJcGWCGH+019QU4l1Synsc39YrpGGPqYDbks8/gEqMkVnkwPh8zaU7tmtJJv6l0vTpCLJFz1Uv
tobPeiQnvIhaCUAkYENOggXBJ3hs587FFJ8fLmqJJCw0sg7drJhLu3wWPBeqzDht/Z1Ol2hyAbf/
0Oq+CVREKY4UbbCLHFn6dT6kirU+zICwU3Oxnni5bOj/NlT+M9OM5d6z3gmusUN2wNuc2FKa5n26
k5W/4VLM/B8WoztDxP9bhoPYDVyiRdtPZlU8TShMFoqILlhDTJHpeVJurGU+OVRjWac7+rNYTwdt
Rp0Z8Md2T/FKGwfX1tnNrq1H5U1vshrx03inmovwN4hEMwJ2VAlkSm4t42awAAWjvGZvpYG1k/3S
4jXy84ZWGtuRxuRszH1B7V0pLZwJ2tCQS6cAOL3mLsy2Y7RNIYI8MNuKG1r8W8PsfnO4t6BsBwkg
aVFph4LT1RprShUgEWH8BBMEg9etvXYZ5Rz+kzZGYF/FhWAijv40DnddouvriUfMe/Y06Jy+EUri
OWAgKJOLB8Bw/lxk0dlVaEqt5CSUN/97+yrnHs8YU3DhqMyK+IVtbsVjwMzG2rMAVwnb0EaAZg7I
h3y3vX5aYw99Zx1AoZuRNK6IGB/RqvY9L9nZOHPUA7PwJfiyaOZ/UGBtkfdqV6KgfgBOp7quTgCn
FLJzzbew908QTlYdDwpsY7BrfWRC51U2/LspDdteBWT4xRSKy90pXXN5nJ39FAVWrxpn4G+ioDzA
mYbcMPoOy601PBmDfxFmrgoKQhRuapedbM8RnkOoibAAPJTEbdMEJkdNf2rPv7zzWsi3JQEqAu7E
X7sVOm0KRJvdgSxcNelKykRInS0jooy+JunoR81CSvrfP7fApDQ8wiwt0eLCKvDw1wlGs3Gj7mQF
dwMBrZuNcHeJc8cuNs/DBOzO+kLDvDw+Pz4WpY61tA3zFXnwy+Gh2VsygdzFoaodXiGVWTgresU0
Gj7CcNnTrvjiUe19sltnC5jF9twXbGbu72pZfyhqXZTOUkcQWayPc9YqMQXIstxJqlL6UvpSwoNE
x+vUSzywdGIVgDoKPs0t1x1J4W4ebKID+sZ6GcqIZuMz1CgMeAPRR6tiH+SJlRex1salZCX61UaK
Q/X1wfQqURfovo/+1c7Xp84OMaEqlPDsJDBAa6rzKphEAdgNweqUmXsxXdwCNvn1+PfyX/lcjQH6
I4JDatowAZl74EOPQjZbaYYbYpBBDwPdkRpVQj8mus6ZSN8cNBmcmnW0pP5p3TUEPuGxDNrzTHTy
Qxxb1Mm0C2bj2oTgZyGmg0ddBcIqm4933HJd3nNgUmBWxnG88RiJI+ZIzpZ37mKWU8t0jA1IbS1N
MvEoEmPLOIG5VHEee99lyV3Y835cORanQE1ODXvosmOWcb/1PVSjBBxF+CQYH3J+fPVTkzQX8NGZ
aRu85sZp6F7TcgvXjuTivuItRXDF9y1Nm11/pg/EH0Kbiu2BsGu4j+l0lXt0b9FHUJNn02LxwQtQ
7rDWxiSOqH6l+Jpnn1DSvvpmsX+dbM8B5qcqwM/tlgAF6iQNzq7i/tBR2zK80l941pp/YZrsS+xn
8Cj8TvUz7GYMt4lq4eMEUMNpZWAueHQIIcbCGfP3Ys6mvPEy2t4/rafpRnKVpx05OdPMBpCMNpUr
Ja6dER4SHnEL+X8HV/45yv42b6toc9XSzPz8ekfdoRatn8Kqei/R1dQ+PjLRsZG3EmJcyjV7IaWo
9UewfFI+RizK9fGiOZ9Z3sBAO3sy52NT5SaK1MlSw0M8oBVV/CPGnmg4MTgxvfrV4acgkfMYphaG
uINf0WA/5zrPQ6QhU2aeOVoVIUuoz5z5cAgVzhpfJYx0cwjcoxWeqj0pbPCwJz4THF0e6TRhrKCd
vXvEIJZUqdscR6suDik67sSDs++YJkaAkbnh+wR/NAUOSfTCMnwjLBiNc2dla5CV9KQdAmDUiW3r
weFS2Z5eJD5GMqGSRY5pphtJgrr6PS8CD3KXGI/wAuhFAj1WXQq/MA4lvh9uwkdy85brR2slzO42
L5NCMEvJopUTAFJWuCXpnx6bY/vDwjbRxule6Soj/7Khq83x6tJ1E2KX92Tv5150uOG6rAuPLpiJ
fFv/Vv4B+BCrlNLmBXgSqcP6zO5NZ4kfiytLL6bnlDHGj5eVlimXFMWGPv4FwH0XyOoLZTYMFH6W
afA47oXpu26bV/Zpx8dqisslv+UeZKP9p5GMTd/AcW4k8X0/aX6Dxy/i9UCw8OFwhWIBjMZ/Tg90
Q1qiRdV1xWZzpDFqvGWouhucuqYDyyibdXD+rpq0cNwZK82QeDPhy+TcsOERaZY9PVsTnP6i5vE9
QPLT1AGFTvfL2nbMHtsgqy1aVQPGqxuGrKKAL8ZnosGo/4rujpepOGhIACTvx3wuyjnzT7/i9n5J
Q1jGqalC+X2B9mZ8R474HZmdg2wfNzkD1bP4cleEq0h1yIZyKFLetA5yUCm3UWg2ZxMDYXeoqfAA
48ClAKC5euF0hJRKKXgSf/++CzP/KAmHsn2ODLiunJli+Zu+KzN4tsfOFk4sTO9wlj0iMK/K0sd7
ORSLw3aWNTm0mpCgjYZCxUh2MZlvawAhWIMIRlYzH0evoK2QnAMnkM1pbHBpsgZsltq+NjKRaXZb
2Wm9Mg11lRj5n72spkMCiCD+slK7CEoewF1xwYLGuH/ILk3YuzlH9qgnb8p6hB5OW07IPV9BJ7KK
ZA2U+quBUnw3PMBJUw26A98j8phWky/GlpmT2Iuqey86iX30k/tS+F2QPbjtmHGb7s6YYwfBBabA
uv+XtB1NGS9MyF6mg0j4P2XMPfkO3dXQPwuyjw7esr5GdA8R+4sGNGzJdYLdJcoFvXNSF0DMIkZz
6wFolzfbw2PPhNNEUisOB4/Mm/XcsiuxznTF6QJz+uuyNGW6wGhxMiWlnXYiRyhqjvIVA3qyEfTU
GwXSXE9UEaMACFfddlB/ag3yrxNS/EbFdYR1dRheqT0hQdBcVqJXt2EGjH26YEC+JQc5Ylm1d1Xr
fC9cDvvi7KL9sTJJn1cKYi0bA2McUB35pLsxM3KmuDTDUFYr770lwo5ooTvu0KS25V5ndFeRiU9p
YRdalr9OWcMS0/4zvE+oSFnAWA04c5r+L4iWYLzcFGK0MON8lUztrArJlBTwjt+ngxIAbqg7b43K
SXAJC8qiyg1Q3N1FqwTtII1VyHPSGQFv0PUf2RWgvi7I09Zcm1Ae99donz0or6F3r/xjdwhL5RKW
AJ3l5hhQgUnNm16wUeIIDtxooCM0Y0K1shMTPtZnnnN7O+KzsTZDUplvnEtsHUhhZhwh1SM9vVfD
kFex2dGER9sI4OTZEgs90vGWVrnMJjw781FvVWFFIPXry36Z9/aj5GL5sc/bDi5hYqR9vPmyovj2
LTfdFumbn1I+i5W4lWGUTpPd/g32h4E+FsbmnmoHFG5i8Z/v55SGNrTpL5HY847X0NB8Qu2iAeVC
RTSm5oqbo+rbqqyRg9Vl0Yx029XQQlwcHzidSn4WVqmO2tB8RD35cz6to6ck6AKqqxuWwey2tSa2
kfS4hH350pUDqcBGzsNuWyUYbgWMyjs/dewjpgXkUQrybSnCbfuVy34BHfMuyd2H81ScB7zwJB3W
0eyrNgz1iBtEL/6BfcQM1d7a2ccMrJEWMxOKmndVqKqSs2l6+xc8rR+xXdk+BduFQMfln83QhieG
k3hVB+Qbyt/tWcq1OetEuHMwsWqTmbrTvk6TfEfygh/1fIiglRObArhm6xi9LBUHsrh0F/xOp8a4
dYuNhgE/lf0ZrsGHZ0vXIZQfoELO23KXCJcDUr+AADvxhKByxgYUQBokjlZDMf60BW/Vz7I3UJY4
feO43WB7o3ZSy4RV92d3hAAzYCQq3VvuEEBLQS/p1nusaU0S7p6WX8WXbvoXgImjhFU1kUdp1n86
BXs7qHawVdROkmWNPsXjFJ0VHxQcZE3LXq+q+NCTaSi7ECi9ba6iEQ8/M79Fax+Ba4fugHMvTbwE
mYXi6zMhD3Dwkn/urUXjwImlURGx8FQayTdyCdCfXUmnqRW4mce/cArIxYvW0kj9T4uplra8hluI
YFFlBg+4Ll3NXuKqvDzylUWoWXidKF8mJ6Uwb7vqMd9z0pEHSi9KWOmSL+z3+BcCfEfwf8oi821j
EcWolu3WO+iMj3u+jOTUyFgW0mgDxUxT/DG4cNB/qdfIC4Ipoqk5NAuPe6UYR3MBNEtjtp47nyeP
1G4VuwhqMZMldv15aKdzSgO0VKpD1bWJRHsZDVd/iNaoBxO2/skdazcYCkCShdTjXW6VCTmjsd9X
TiXgGUlRTa5/AeU5K9rEd0bc1x813ankUo3QJqGWLlp9z7bFLI3AQeJ9WBlv527F8qXAFhcYAELw
6W5CpDAuv454Ckfk0pzFYAAO5lf/SiY0pTkfPTyntRW/5AhMwByQLY/knai3ijQjjt4LFtlAj6dT
YkTnCgKmxecppfYzqLq/q09b2oq5novOJiQvsUEsqxB1A8oXGoFOq2ghFR9D7tyTfI6nc24UPwQe
ubZjE3CwFyv3lhoIhZU/KCmuBFgnFLMdl3hvYNzWX9XRVC1XzbRagmw272373sf9OXyND1U8ZXJM
XDfWRwMoFpW2o2OcWHYaADp2eGfOpKaAgKJMVMNhMduO7+TZyZXTkrBUt7L+WnTkMUHuNOxgfz0I
Pje77QDaBjsk6i5RuT1haOF5n4c19QjmgdrVWjwqQTHttfs9ZIgYTOc8kXn/vLeX36ehIt/LRM+7
gbpcB7w8+yHYsVkW1DewCrgZXBq8AV21stu6C2Adgu5zvNG0q/gmWk8Q8z8vIpjjj58f8Hd01LEc
3I+4jQVRPDxVy9i03ucjnAz8M3q3bx/Bl3cQ9MbtnY5HZ6Eg08FxWvISnM8YlA8stoQNIz6bOZbY
OJirkayBowufPN4gtZMl0l5LxLIAOX05ne586UYanZRaCc5kiq8Q2vV3yy/9FjfgHzuaE1h0bik7
lXOGwtkMXR6EqI6Cc0GehRKHVL9ppwgBXEwQPGul5RQo+H0K1JFWKfF1x5JnQMRCh0TyGbeX/FBa
3/QEwOF5uHTY9JTAvpV01V90YhM8UtgLQqZqWdGtiAKkBb5JfQ2kWLi5YlmIcmXNVEd0w8y3N5QJ
kSSVbWRt4eusO2UeFiMni13PlJ7DGfgE93K0gSKfDv5R1rls3fEyDM2Glpu8UBJD+aZwEMlQf7V9
wv6n80lfu2J9c/4Ps0aZDtOzzPZtcnjwOerSPl8uWKNI9ztzJWenjK6RVvIw1CMN9JqaPaZxB4kH
otjA9cATIqL52208O40eSSU1zw875ImIwnhXLkv4JFwN1+myt6H2Lrg8RYJpCV13CTWPYwLeOMg3
1oQlx7JZkBQSsZW2Eaje3RcVkPMuhs0GI9XekmfcpHJO8QeYbcokVJVAIqTk96Tpweef1ggccjSE
z6Zav2CUD+qrgfST400p2sfsNHNGssrPp4WcWbht/SLv0AS4SV7bd6cMYFCj9v3rg+PtjBxrNuRt
bNqcRWEjFzi8YeZ1e+gPEVYlccDHiHPNwO6WR75W/dOEtVcILadPyRDtjVG1UZAAomFnBLSe5YHC
PJ+fabNAuE2l9Myp0vaUHAE2snYla3vcdP4fWG5oEjWNtJ3aZ4gOe3ydeABXJE75Lb2PyswcBZv3
g9KoMJmVbHNRGuG0TitNSUDx9W6v1T+VndkeKxOAPwRJIWQ7eftAI7apKxnPAjHuV53bqcdXkEXm
pzWyECDW1/zZ82ndUdMdWXq6FzNzGCu97hkVry5nUnZSenoa5/5zgE0SOHEcWW7sB695W/UhbKIr
/+UxYUDXADMo3O5i+o3OIh3IqkNst36tRyqA6+qs0WHeQYbfbnbtDDiMxifA1rDas+Y8LvDIKhv5
obNwpWlIu9cuGfwnT0sAnu4Xv/s7CXZc6F5QVkh/VELmNeqKRHVFoNdfe7cq1z4EmxFFfU1Blsja
ZOE65lbWFmmLM3igjKX6JC9WX6UUdX0qyBfU9LTaBFD2YnOnHrhnXvmA+94wGDLGQa2UEMv3OoOC
6TIVj16w23uDde5WxJN+y5AUJOXC5TMTzEB7h5p2W8pVexXKY16zYIkWCmOoO7KtBuTNnoOlEwmq
4yHiy2oDkTpnWdsiYEKVnLFHpm033T6/e2jB8sYRgp7+rxiu+TVDQQyqckOIMFst/Hl4T6+0krs3
sZH6YtC8iagaNn+10Ttn+kWDxh8xTofok/AAdMAuRrNbfrtLKHw7MIfroXdcoOuvFin+MzytF7CW
ctpNX+bbgTojhpGEGl5C+greCb91leLI6v+22S6jYV9FsL021ElbJ5kDm0PYXd2Zf8hSoLfvFuRj
UHLFbHRuvsndG9qbcWxlAckBvF7L6v29jfAd2pwS9XvF2zrrBgtoaTON/WQG6rWHkhg7JQa+v7lY
B1TF9tMoZTD1o0xyuCPaAd0yrev4HsNiK8iyLbTNt6I4Lc8Q3v7I5kwOpxgAoMO8UqWacqlMnoWR
PAfJGNg+NC354XdyG8cQgmoWMZpbmonRThDXeqSsdQwUEy8e5zMqoj5KrPGNWJFtZBTN9jgVw/wA
ljF7/CK+YLw+gclAdao0x7u8xyLYYiBy69OS8e1y/fj/enrpQjq9VLhtI+xKj9OITgTDrMeY2AJV
Uy+9pQXUuq3OiCzBaxZmgQsHsmMNKB4yxrZ4KyMrHGJPC+5qLzsIPwFLAMF/9+10L56Q4yc1E/NY
TLEJUyLCbTkRKYc0B4t5aT7DBtiXnOURnacL0Q5gpc9/AsGt2Zazj6+kk5E3yv1LvLtN1sX7iN5P
P8oNO7w7f1rkked8ZBy7N3bq7J4qZd19CHlBwC8lApgFNM0JCxwRE6fmAqVV5RdH7g7Te/58xL4y
V6iB5ko1VcVZmn6+l1+xvx52q5DZZRFXVCjye96T9BB214WDm3/Pu83EBVbJZz6nIXz/nY789yP8
IdxLD3ldJxvuMjNgpa6lnVVxQEPLcQvWxb7/Np6HitInHAtAFZRQMi/6FFokWFh28Zl7rZMaiikC
vhM5mGGvyYtrMPd6AkbOaaxkt/v5qCcYVxuclG5i6zazNRV8dYcZRgaPf6OOgUu+srqs9V4ll22v
7Yrw3P4THCZmb9Cb2lqUwfNoGa4WgJ83rDKPthxpFXwXYjxju66s4hrLMlyGuXyQIkUhyqSLGQw7
CZILrIpsmQhiFlxGxcGS/AzttP8W6m8FsxRfHGallAbFK4BdNBw1FsIWjDgOuOF3DFs1p0HhflOK
GDE6SPn79tO/xY4hygDB8TvBZoQ9ZI4z4YXOynF2B93XGO2IduWoUtIOSytn+u+2KP4NkkQ+xX6j
TdExH2LX1wUSs/3vAEx+cr7wjBQz3Pg72kMuuGX9KMD1a9NBsMNtqgnR19I9zvDGYeFVQoLLBBcH
dbXFl2DrLyw5X3AOid5/ErwAsLV5W8B/Rd2/SjVZrnLt/hTG9JzPw0kqXYmEjQIYLDqVUKYNS69N
JoXmBBLCu/NBK30w5WLhzIYu9JRCUHB24O0YyRLCUNDqG/JRUUgjOxle0LGT3qdK1hfYRIQsz0wa
o1K929xJaPAkeZr3Rai0w2TlkVXbfJPOAC7peSz9igPr+d9K2yY3HdoTqzQxhyyPBFtqOOzYEJ3i
sVGJLoGSMYiTLhMFdcYOK2RxcJCYgmKGb1oIe/brRJy9Qds7rIwUGnocMgArDuPey0FssujxTQsa
JfWAQN92DqNsIgxxmubHPFz45anhEgqIHUvwOkkqt40qogK+s8NINZ8I7waj4HgmWm6EX/hFI1Mo
keLxLjt7HMZxbIgxphXKCgEJxgSXKwlUPHzx2yhDNPxSG7VJou7PcwSq7fwYfuUpJAQoi8v85Xo0
9xTXpinVgFuOWuVT5ZVLXZ+6SfVNUiN8T4xKcX9BYTXk4KkQlwEqqXctfrmzs8MaAuwlbhsXfEY2
pbrsyS7qnPx4ZqSvEelTkCebAnKYywqwe//FaGkBzGm/Ic+uLnbOdARjGn2jBE4SbXzC0vaCKxKJ
L+/MWaCWuvvAjT0FyMTOJE6JrqPvLFwco9K0fv/84dM+W89HZJrdw/PVZfFI7+o/gVIkNZlMFz4j
S9qhv5qeszglQs0g0dNn1F9BkEJ/zh6YGafCBNXayP3GNehyYYHrTp4FQlPpGgUWdaWvtWkXTkql
7r4IuLGedK7eIi1abbH0hDNtzdm4lR9UY4StB5NXcTrpQVrTpNUN2bD+iiTh4bjMj6zEa5MV/SgE
JbysL3z7dOVQetaU9h+Po1iwLB/HTPHUd5os76Y9cd2jrUXwwzIvEZK4VFb0Hgt17ipYZZsuVxzn
4cVVExy7X3NYjqT1idBCsK0RMFVGtzdmew92SmZ76Ywc/QbmCwBfqn6es2sCcE4J2VmyGUHdwfy7
+Vnk11pY9DKuZuswujU4g6GZN8H6ZJ20v93YC92qp0pzkTa2RKhGjmLGc//SqWZ45ZHVHblToT97
EXteoKx6sTVAWrtC5WP7ig0y9u1Aq2bXN0uAPO9prwm9D9kaNlgqk+7mhghD8ZrHKBSyf+TLfbwD
BWyoEhHyw5YMzmJMVjYAwD0LRtAMef4pbOCbsCfWpZ2YEdYjdObDHa2AjLi+DCGXfPXi562KvTlk
GK3/t6JCBADLDqJ4ahgIgJ567JO5iW3VNor4DYaFcK9SCnr/X+D34rnaB3MsBJ7988j3M5MNxBE6
7QbrLyAZVc7bLfwHcDWGPVp91u0ZVMANI26Z/z43hLQZbKUc9UNFmMYp9QVweQDy7QxAXwReNgEK
1AwOyVB4hbd+Fl2chjTEfXCc6a+/fJYpKkHwoX4ZGJ4VMfZCt/4AF9c9RwiQ83x/wB0GRBCe2HDF
YMmgNIShsAYRl6wX9WeC3zTslOexRgSXZwwBMv5cX3Q6Y4Z9BZIM5LTyT4D5t1VsyBKw/VIjKmK2
I8BxB2klyzXADjz0KgN1DIx25bhKzo+Mjsck8Gbu/MKf++4thSlpcrJNX1BHNMJESBM2PObOc94I
UHgMsRdXOcS9I4gaU7vnqsvcae1CV8gjWU1lbNxP1LYi+luKvbuQ4fLXTlPVS696eIxgROsPzNV1
g+dX1Y8tgqVDOrRgrqkzAINa1hUt0bQpBgGtji7NJkqwcWzWtkWgW9/Rs/TIlDDIPRK9vMrfi8l6
V/7IjdpSLVIK0LnBAq3OWbhKCOCNKNK9AHbEJf8GxmszPKfUXjcsq8o8rxa5AAVYE47dhVIBZir+
ARITjDc5+uZTXvrqYTgtTE5GUuizYAf/GU7KAM/kkPoDIhoWBk4HRJg3Xl9IXmhKHKvh4X6JGN1n
hQb3ZSN8uzslz1tZkxGD6uJSa4ul9jHQaIGGNSS5wIxhj+wSesKbylXa45GTSJyhxrpkcXaestBE
vp5+QIB+uvNNXptkcMr+pIIwPwBzy1O6PYc7/0CU2TlvN+eP5Wv2Cxyhb5jpkZVwZ2ftMRhrSMck
UzY9gx0G+2RjGkyTtZ3GnLn0L1d9MDEGeoR8ugcGKFFUz7vAgHyUwjWjcy3U0bSwFgjCm1o7Hrn1
8CLutUaaP2NG8kbKmeZvjG6ZpuTVxWRMJoSSsFhqbthNboXYLT0wD7aE5V7YOIXJL9qxZvRCns4Q
86pQE9bQZs6MD605+049pWTdo+4BSlr1fesgQHs7+wphJlcXT6HHxepjo8IoUITRlq2rIWFP98CC
g+loHo0w3aNjM69qSVdnycrJlpZMImHdipngxr5eelhJu8MGclugmCzO048sKpunGx5gO7e0RH7R
7I+FezBSa1xzHY3J2yqpG4NYIBiBpywf3R4q99MU76F2XO+mjOrGKeedqXjlqTM9N2pZ/r1wm9Li
W+kk9sJHm9/wmzA6tv2JzZw1/M5OhcqUJO7HS7hD26K26k9qbOy96Zh5RKZ9TB2UEvnzOac/sid5
CCV8WS4Ko4AWBoAkaDA46K73ILK3Wwop38xDWSNOWYgkxSTCzwXZI5V6u2UkfOWeZd1oXj7jDjjS
FGIE0pwAlCLwocbiK7mSU/xL1hx6FGOv+lQWYvQkhBm5tFej7NSAmdKqCO1IRQj3Zn1vXLAbL9SW
vA6USSrICB2uLEBQG6B/Mk88WUHhqeGSMhkX8iTKCmh35c9/sMDcFR0wbxeuQFvTZdxTsKJl+1f5
LgaNRS6VfPtFwP55xxNK3yamze86rIzMUZBo8dMbDDXWyPzd1L+ykgwfSaFKQONkxWHKfiz+BeV/
3ro1k7MzCtEo3nhaYd9XemxobWipvM+bKIX+AzzaofJRg2CbOBHv9a8KHZjkJLOzHSUSAlcC5WZ0
v+jvrBY0FAab1ukAVj1Az3X3R3t9IoFoAdobdjA8wUgynSBRSqng6gkit9jX3O/RqO2sFcF13HNk
Oonf/cCZ+yIzVwh+/wJEwH4jqChGwL6WHQMvhDAheEqNCGi5CWJDPfbyGI9vaCGIRWVeg5e2gyHo
lZSbW1CD5dtXYZwYGHBGUsHbyVgnzgLOo/aB0CkB9hkTOqORp6nP21ycDk34WYldYR5U0LzGCy7K
vGRfXcgN2mFKyzV9360893BnBJLd35e61dgG+Ng3qWTmyF5Qr1kKXLOHm0eCpOQvcqI8hAIH8gRa
KrNnbKGXxyyv2sOVJn5pXSV/JBPU2tINdLritWqGPvGfAp8NROQ+sk+TFju9wSt2UEYWjaPMYNC6
xLJFqgSxnB3uVFVaGwp1UIWoa66rhFXJ7JYnvonpq9ONjyNxR7URXzzWobn8p/YAEpjDlD8sget4
DqplSESGs6C807VxBIt5PVObyXij+wMmlYHPhCb1j+tuIthN4a0KLy/pZNyhONKMaOCArPkUw19+
4OsakmxG7QtSPtsW8kWUIZuE2+eOj3Dth0k3nWOcU8kez/RNcYsNlGMfRTVaxMtn9amFClvxS7jq
sVHTGyLA1+t3M9ORNjOt8uX4dZClDRidQN4MGMD7SQoi6vF+xKmjYjBL4Fh01HG7TdaXdkPb0OfK
7jeKmtvpiY0j8q1ScORJkC869UvnexCOnysN4LJQFKGwEfB38n0+ERM/pHIbSZkVVmMfluUmX011
0gZ18rJYsn5+9bVelBVtYkyyh+s5ac3X8QfOtj583FOk2bpSKdgjBKv3gyZjpIvcAOrCDIJukVT5
lBjM/EHcoHIzEac6r13jYQxkVuUqSlzhNa97PV7k4zgAt9Sk9XSWwHV3rf+Z51fpNLhEHYVq6lWG
Fj2NBY5mtQPyDXIi418gEY3I4JN3NzU7tAuzkWUrViLxPoAZ/+kIAdtWwaW26rEvEvB5Zrj3mPAg
j2Qwu5kD+kO3BwkMhzb7MtSIOS3aeC7jvDrUr/Tsv2ze8kUezoM3pb1cYFe9XeH7Tpjiw7Zh7qIe
qnudBPOpVsqjg2q2Q/8/JnBwa2JGYHM1PYxEDZZIuTe3czOmslpMGS31AmFFSaBzuRtkYJ4bcuF2
k/EZfiSFshxyP9Fvca/m5GpXh2j0CjebDlB4Hb5HYF1mk4gjMqrkIuD9OzFRv8aFv3ptKHWWZmRJ
RbBB1gKEtLH+ywh3rvz9yxxb9CklP6Q3TFn0QnAhE0e+qLEaJKk4BxVDQpOVAs5v69PhVk/l5vAn
vvhKGdkXSUzT6zwmBWKbIt6eTxIEQoYIHt+Bp+6CbCPzcQij6oAGVWNuczTDmkAMCib0d0bQMV3B
M8lsSPpN8xqhJQPGrHC29ucyfiYxtDMmKtfccSp3b2IeALoMtkKAxug10IMQtgJ9DSl9eBnQin64
tSNa7IXnnQwQmPSebD1LVALmx52epkNyV3b+3/chMH74MvWUB9G/rKO1YV0WP12LaVwJLPCFOmN4
keNztvVjxHjA8BK+xR6LczS17c4cclHCtjkdP0cB/t9XTt0V8eJsjUZhThxxst0yO8UPkVHCOIOr
rbgslpLsaFSFOJHZBFx3Bm70yUisjn2YF0rKXlq1k6nIVshtdAp82aqFaOCuBmsDK/Y8jTiwCNfx
7iGWZvdXxkHV+P6QPzZQAvZZxnwHG65Rq+T9vDoCVFjwFgMzpg9e9gBc1fZNyoVnUXoKOJPXRmDQ
NWquvqiImHpCwwBxHpGd9KpyUcEVw/7yIEN9XU0LQcXYT+f8np12mHovgkbpqwNa/oYdge9gArHc
AwKxjtP87QChahYxKT94SDKmlke4Q+RswiMn84J45Xv7uXsA+til+lhFblc3ymuLKNaftszortST
4cxW0g446bbroMzDhEXn6H1yxyvlZ/+yt3mLyrh7aLVIM1v91FWPFs6PbtjAKw3TxsETxUSvfLNR
xMLkUVd0V9DOOnAeq3QYMcGjrm9qgrkIIzPKnN2rpBKkfNy2Z4Fl80habO7uq+5nARIGcyADgSGm
dMFIjleyBciwsp2AADZB97nsFSDTJ7aUjTonpjusnxSo+9EWLie7baa4medB5cQGVweUjCZkB0WH
kpPUNprDHnNPqOxMxxaQOV9LCynQQ9n3o7523ig5OVOk1E/eq6XP/ycVF/tk74QtNb5kEkhJWNWI
Y3pTXk/NX/0tEjE+p4T3T+ygKr6q6ACB+0jIj5Ca6R8supN4AXhuhFJy0ecE1qJNvTMTwwkqx/S/
riC5fjiv6P8pvkC4owrGfhaooJwnZ0T7acUBago9XnX/wZc2KhFYKWoyEDYYhMclbObEfg/SjF3V
pgaC15IDBbmtOhB7VF4RhC8aey3gD70vukGQE3HvnWSXpd/cMBWO6VMS4aK4qJi79W5e41xagyk3
7LwX8RAWAmJEEaezYY7dOo8SrTRuy3PgykAhIqOO43m1u3ZkAaEHwbdsMUYpMduv5NjWoJvSBFkr
M+U0S4J95muwcIbV2jW7JD09NHo3voXm/vmqAUjYaxDsSuDAt3e73JqI2R0oh5+rVK+T8SMKmaFn
8e3WBIS2j903jvP/ucLPQQdLCQxwo3qkr+XzroH20RUD6aubO8WIM1rWofTi0254ucDij3BE+1Ic
tE4G0rrHBDfCWNbEn3BWdo95bV645QteAygnWaJ3dZ0bigOL7loAC2m0C3JxEgMEJBWFWsEVZI2W
cEFKSbhhcQKvqDXQpBtLthvscmwWy3L8pPCLQetykGvsCFxmTziVMF0KFYAX4OhbCE6DCwKr1grQ
pIRj2Xcsdw8guDnTHkocmO1W6aEHBlKCBprfei7ZZ4Is7r2GBF87CGxX22mKI1JP0ODhOxH2IozX
AY+/gTDX1oN0TCgipHEI+tkufiPImdLFOtHWKhGge5/04zffkS2JXPm0tf/C+aiPaF2IS1wi6My3
4LxTKgbBS/JEkipD825Gx8qj7DISEaMb02gCW6wtnBd1TEPgBLmBS88D5DtX65ifcinUpaOvvDem
b1/GVGrZVwUdP9KpMZaJiByOdrGE4NDpFU7dfusFIgD9lX1wj4X6QTAwVuYMYctHNJtHfr5/whQh
5GFD+KmFYT/LqWruVB7EECEe2Cos3k8v6UYAy/zXCJr7wbaHBZRVdkWzCJdShbR9E6Pakx37qHob
iMochuMjZXLxbJ4TzVRzDiG+OleGRczGorbhesLBUHLpvuBfAQ7zGtkp1GhcXtFn8YLI4uIqtezc
RLh85DZdnpLpLg4qGmnoHiBfbastQ+OhRvwIrut41WPTNOMn9LQCwWnZNSdjoeorj1FvGN9PVwrb
Lzyv+UgccvsCyZ7GOTV+n0cLpsQBs5+sfLJmxYmiIMf7G56odjOaNnu5793u6J+jNmXJFpcoHRj8
RzkWFeGnFc315nc64RdZYWFB5nsP6yO0ZYz62B0ZFp6Vw8cIrNYqFptTGTt+lqfN696I6ov34qa1
Vqhi40kBy/4avH08zchzn2F7BSyjxoWbSLziSuy1dL1TMLHhSyGlk39jfc3KAhG5odZurC/LbBB3
T3V0lLSOfr0it1T5PzhSPuznk95vgw3GEhrViRKoa2uYc/mRYPha2vGt0+S1idSdy5JLNkKzw++A
ksUlo8OtWS8GQeX5VU8TfNO63xriXVw2e2foRyej8tgIetU9BdlwDZM796WApCe/N7SwvPZNRP3t
EY0lXCPsXdvCS2LkPNft/JdImDVhHWDG2eVacVRkcJSGJHORA+TcOOS4e9M0s+kKU7DKzgsV3Per
jAouLjcDYi9oCdJOfCgfUQlu9Ko/OPIWRYOH5+g+Rj2g+VZvALnSlSzJ3v+s26P/fLpRv5YnB9br
KWzOISYzAaJ3o1pnJza3rKps13ymfjnLYGOe1U8b0EPLP4ayYNoqrjds7Eed5zxLWOQjbSH0Nlyf
uwq6NDWIvFPOvkxQf1Ot1vy9ySGdKJQayQPOMtnI4n1EW4SrDiZVIjD+etKTIVHnn7Sg5JnfT/qE
MUXe1qDtqPRyFj36SRpd/xlCSPUWEiShaZbgTD5x6RI+pU4lNDSjqwHmX5IPWIvR/ZSQqZZkXL15
iRhfNlGUEiKw+uWExVpSNYI8WROznSdznaYiTV9D3K/HhathN+XDd50vgJ+qvRBPI8t2a4gin8On
w48UHkrZ5fb+YrttEpLKWprH9FqjxNP4hGMm2XZxh2aAuQMgHHgLOFWucpChbi6pXLhJbMJpaDh2
BA8UeIijbZ/TKDgjeA32gQzXn+QXR/ynxjY5LQbBWDunr/9xfS95ZMkcHxtGw7ZnnXGbPDpP0kn9
8HUluKoH2s3rNfagIiCFl+CQjJieV5kUbu8hA/IwpFM/D2g3ebbF4Xa2uMsjBeU8tsGt3/PZEFKY
0RPbxqeL/oSkj/t+vbfEx1XoRS7lvn/KR7zKWbyUUp2nz0D6jaJY+kIPLn0sBxpACBXCK/+Cr8Yk
wH3P3fMvVZPIDDjIpnDa/e1nmvwTXnHWfjAKmFePDdT4UeE8Y2Dv4Kpr2XZI8PH5ACdLKyUDhC5z
yChNOK49SogAoccLkR2XXH6ONG/WEZH3b1lJWIaiMsvBusXwhQckHeIRzcupXUG3/c0dNdD7Yeel
QZ4V3Hyr5oV+rCALPXJqLl6coJCcwvABmmUh6+0C9L00MvvLVmotskuQLd6ZsmT+etaSmbwtTfZL
XFUTGFspum1GkEUF67iCOtmOZ6AncgKDJuehcGsILdp7tJEpr6lmPTdvQ8eLhJznLTPLC3d2rUZM
oRM47j/XeaEqJr9Trqq8OXe+qSD8i6ja2ZfPvZ3EPewzrAX/hiDqJ13Vfwsc4RsylAp08ykpCPna
L1y93msu8Y/jhmgPlaMzmjRrGOfKr8Ozf1CuydujoLKfFaQm4xLK5Q3i/4EI+YZPPVs96O8cQ4DZ
BPUAHJtKzPLzkJwwMTSGNvB7C3KPRQKL6pN01gOigQr7wSqUAwNHRXb1MplYrvxNYlzM/HkzVmKf
kvW+ajYdMrPT8G2RWgAk1zWbBNS7TUCVZCvdjJg89EOf+15Xm2LJ04xhs4YjkqB3BxOh/g7A3ONj
v11z65+ddzBx8bzpwa7Ae7dN8y78hNZxIW2p/V7iHXSdTGrC5a8n1Q8ikIEMxZIoG3K7lJd0aY39
GAJv9gfQHdQD+ikBm3h0dmBCYvklNAeQpVwdabgSo4OoEPBQsBGd3JHiMXxzLa2QiEyj7LDFT8Ai
R/vfdQV3Hyg0tfDyfQfSBg9mV+NSDKmheoO5ZD19Zt94SDngSRSj3/T/9qLKTVy/gYyYaRC8741C
gHWRBz4PLRqGa7f3S5izCuiDt6ARXOD6ff+D7EJEU6CcIhSwZT3H7JvdSPNaDd4v0oJVNPHO165R
mxKnwrAM/oJU2IZZFarzKTiPL3wycecduWBTnsrYi+jizTsobBTDuizORuUKm4pl0d953B4ex3gK
UOAswtKQOESISjtNPi0il5bhol0cw25g4TZWlfgp42N5tgAY9yolQaCUYkWDoqOfGH+BKKDi5qPm
dGgiCir0AQlARPVRyCzDchKN2VIuEkiTRViA8Do+fWjEmKKUCihxSLrHR8CZgSFrRuICMkCuEK+t
KonwXBYMFdtjwsUcN+5oKqgtnaxB67SNg4UD+BDracVqBfKDRWpBhpAa5JtSkKbguHV+s2+7q8DP
//rl4vkI3nHg92WuXBAtmXDdLcUzq3SaDXaLsvbl39Xdj9w+aq8XKjrgFf2fOauWFYQ8l4zO88YW
o94lErWvBcvj1VqH7psitWrXsIh9NCNw4Cj5onUvCWeYPfCRVmysylpfzFtqEyTHdsZ6btRbQCOH
eT9fLkQeRE3Ipoa/xss4nz39E382uwE5oWLqsJTxPtuWp6U8PdEvKR4ADBX+RjRGEtfs6nFPgk1t
e4ZOyJQFThBTfU+t4WBxbDKwk9C1GOUkN5VDcqgka7UNodr/p4ChkZvUPftb4IZlXOSKk1/L2SLV
KerIYOd5DOUmetI7KMp8Eae9lvN7LfLMQl/OYXbv1O2c1t/PF9mg/FtYtLSBfq5tfO0KMmkDaLzk
rCM9QUhrFRNxts87fRTKKusyte3JnFaZtcdMm8/AUlnJm6lrgNLfHB09sLlMf+zZDQtHP2DH3vis
ppv+fhJkZAaZb6SIbK4cti3oI9yw6S1iryyjwaNBFfZs+Cml+z1fTEkihLQwc+5Ytp897c76r7KG
D1gzVKGMqUzzzqUWCQow0uHlphtwkwr0YvsQOwpJtOXzpiwYcucyKPCmNbNFvto/T88jkyEmpvmC
PKJI+/OAW6heQA1heOfdSQ4CzOzBA+UtRhtB58xBaFQHHcrp7btzpnS5ozwDUZDIp/PRU9fiYylu
7wLFaC2/Lx04IEX0hPqhITRNiNQzZr6j6mY/wqMd2IlDdjhv+EX26whg1Gzu4WhjZFH25UFhlPA0
SLMn5zIvPJnfG7PPzHorwM/so72W5tvPoH3TDULRpMJLu+0+Mnm+X5cI2WaxqQukM1D0qUHE9vRk
MOHSDzK5lgVQ+tb++PWRx3IdJj570OHnn4iE8DvaiAPXTc6iW8cI9Cqf7hWha81Jc6wkk1mkUu7x
1oLn4OTcMYDXZPzLAOEg2gqscgqF2bT0N+DNjBldAbYr09x3xufLlq1VRKT73zu+uOEjz92tzlRr
2tDOBZQLQL7DCv10/Btc2siGCI/IXzvXNDUYZZyDFBt0oWY6/6j441WupWF2L4H7/noSXNNEHKCH
yA1+summC48+ClyZzrGZlOuvQZo7IylzIKK9wRSTVXKkbuSuvYdG7iv2iyXRkmW1RaAqaqLgJ/1+
K4YnqJUMq4vM5P7MKCEPc2Ms8DcuT5B8p9OJI7YMSZIu414tr779RJtzDPYwUHwGAq1ICnVfZx4K
tgfI1FYfguZpZOO9SP5ayIY3n2G7Z7ulcqxNEqf9h85b+kW/3rLCVo+Ga4ojGHewVwIIIRQIP2O0
ancTVpTeDY/WbDaYKaYMmIv2jqaxmTewTuP01/SwNP3xTVNPc/CQhlwJtWkdv+sR9IzsmXKiPunu
crGI6W6X35QhHIwbwcBWM1tVgcOM1Ubf41dW/W01Fk0IkkbPg036rSiUWlCFWd5N5jjlN0UT7Y3V
fMz7AT9Zz8LZ4f37ysFuSWnZL7stG8UqAZFPiWaTxDXbSBBfxbinc3DEncVDFJRifa5uDNngiI1w
ND9y7E8ymMyrE84Tx3ELIPxcIN+gVRY0GrNAK8vCDTRMmTsyCHRZ4i/8j0PQY3w+JrQTDBSxd8S/
LtEYMYckS+ABMi/0TN/Gqquh95NgseKXkox7RRplJD6b/Hf9e5kxsqe8BgmZkuJXzmuWHfFmwDCz
uE9Aadil1hEeL6kKwpRLg/kPVCDlyXlBGsJxpWIMxKuwp74l/k2UEpV9nDdq7hGVmsv2PbpwWZxM
Qrj/W8V5le4N/GmxjAUPWvQi3BEw9iPljERFrrr0LUPAu8l9Yo7/ShVDosNyxLrUZtk5YH5daxvt
O9fCvlAL8reWf+EMK2nunN53CV+gTnNqHbKqbhMsD2P9sP4lhjRpEqqZ+Q44Afv2hhwvYvHeoKNE
uCIN+CdRjqPNNZjxAEs9lTujn1tfDd4lZdVDYBGcydvV8sKYnsiEJwzqBTATbE+0h8WkVkMAhTVB
o6pSiHt9BHQpTQkNSwv48Hvx61Jfo7Cf2Tm43EXiX+5HAbE+icipHywp4XsNxETh0jg4sEA8BBpC
ZJtz94NDQ9XlCQOY4RRbjoSATTgdkNyqJltpCsXVJlyW8zlUBXgmZFEzc9vKVfCpIQ79F0O+s+zz
9uyEBAG0CFxyC+qNS/jR3fj2VPQMHruEDcCvtzsiHYZIJtvNY+ELubdcypehpgJ4MzeBQFjSW1tr
7A5zxnocsKXvjiP4dCSeB7XBvQYozO6/niz1ImJPTGcZxNru4SpqM+iUMdsAquIoRbxgQ/oTvhpx
c7eZ2wPMxrHXvDhd8H1nbYXh7txq+NrtLbsxfkMWDo613oIFR0gICm2cgRsgdgMyLDrdDbpGoJb8
ntYpSKimI4fD+mSzEpyjPCZurth9cNAvV+TvbrjRHB3LQxFRlyPiHblFK0tz+JMdXR9uU4SMwWWX
tkhxlGOsTDfsSfVIiRaOq2UsZC9XRIzmA8nwZmECgaQu1zieMX9B/+HwMh5QhaDhxMcJfjPh5VcY
WGfUxcU4vvGcRO0CTQkl6g0nPbIRr1M7GILWfcL+BSIT1xTtwLwtI7v+BSbhR0lzvEl9hHTRUw7v
hxzOA8684Dcy5Z3KfD94cgWwzqH1Y6sTkO7AWjs688pJfbl6ir89aSXkuifeJahX2A9ifBgBszxy
PshwE7i22RmvIPwiegy8KacXourNRUyvU0gaS+zxhNkt3aRnBf22PrPHKlfZEEko/22hCh38RYjU
7/NiHU1zKFb8LHkCyKm5j8G4dNTI4Lo0j0ZUzrlT0zWSGN0UffhBKDQNIsAZaAPiFY5vbYalfPxn
Asg0nIaHeTMph/nhL01Fk6qMQNEw4bcq9eEnY/Kb7QhuZB7zy2LtLSeueH6BPy3eDIebK0apo00n
5Pfku5OZOCXmca5IAV07xOFEMmimpKCN0SQsKHDkhqsT0Ngt03CbbXM6GcZJjkybG6x4Db6rocBE
bENEVD9PCHxGzHbEiIY7NziSF4ltMJKLBIrfzMacRcy5C8xevHdPC8pjum0gE+muVh7J/z6wxcpe
L8zjeEHngqCXYY9cXsKUkb71q+uwt2DjtFlum1DITi1LELHqBynUnOhhYq5Qq4hyg/eBCVOcG3yl
uwck0zHPt8ex3c2f9UrCg75L1kbt6PnKg/LNpFR5csh/awEXTX9LcEq0J8k4lOEVM2vwIgs+gphZ
1kv1zw+XmlGPjboWgEjGUwA7uGanrHj/2Hiagq1wcCDedHqdJegm33ls+sMfW5SnK20aWxwQaPiV
sISXvPEzJEAK3EiohRufaZQQK+BvkT4O1QMoQSEh3/7i35ewA20UX8ShSuyD5zkY3zhAeg30yd+p
JqHIYrIT0zBYCLtSZ9P4A+ADWB5tp08EhfhEJjCBj2kiiu3qfVPKVTZkg5hdvai1ncYerintnJfF
9kdUpeW9A9ihR1zG4BqQ7KnL8yjL8RZDw9/IuQ/mIX/jCrclA17Ccwh12tp1TXAn3Y9hJWUJ6wff
qY1d43ikaq0JgyIBERLdREjwE8gcgJTmhZy2I4aRowGjlQucnJFniokj8GTKGOTySLmCtVaOGqPa
jUaFLeLQP/P1hXNHg+LBEmpiMHN2efaDMWkS6RFMXaDLQPBNX+wyXp5JtoudAhB8jN90z5TWJBkQ
lQQbtL7N5Pl1AK3faKvXM6Mdft9J4/1qN42YlXOx64ThS2yCMI04RM+I+ioiY/QGM4lnu6hgRKNu
ZG2pfA0PSVRRqXGJ5EK0h3LeE6qWyR3xMKl8XQNepPQXouHv3I/dUp+534dTquTqZbc7NeY/i4hE
Bt/TIl4Gdw/dCMGiAhaerQoVdAoXs0J06i9BSFpYlKPF2ad4FcYYq3Q4KKo5iUWWCCWwO+88b49m
h8SkwrJVriCnodtlLSrX0h8mIfXGN9cS7LMZHmh2erXJtUL2wT+WYgkE8t/1dxRAHe5xz77YzyK+
KmiOq5Znstj02zTqg6L5SVmVjFPf3oFQtf9vy2ptZyy73E1Pu78rjo7r3NoqbxggQn1fPSs1+/DX
XxvUAdiiT6RLMSPcTMJbcWOefyUSLhHEDmOXgUEDsHs6T3NTvINncnrse2apsZ6qKft0djZtpNHV
ivieV4FsVwMod/S5g9TQhgNE+4G2pDVYjW/IUewmeLIFa9SzscvpCA2tkn2glJH1jROERD2HX4E4
zo4Ak5llU/f1y5SSvIF/XSfB33dTw9uDAuReXU0cz62MZK44WgekTwxF+4Egu/iCLXVQRaD4DS11
kuNG1g+9PbaiECvLFS/9c89twZRu2qXg7oUUjF6VyN0fRpQp/J8oDi3jDyUh3XRrKmXOnkLYFT02
c4MoLEIsTVgV9+EFqHVDIHRElUwSgVPeL0OsNm8zVCkQ1IFGtDBJ0J88EMUVgwD0Us/n9xzFSfXM
PLFjAm4StU4Q4RkH3wgDS58oUCYfwzes29KZO1LTGybpRFMrLkb2J/HVRXKbs9s1cjGMjFS3J+0r
ZouCpF2M6UCIZd93T87q5S3nXv3CVhy+amL/esjW4pJQHG6yVQJRxXdYKuDoQn1wlaI1PqlAmm2+
im5f7ebGQ4mbWy+/9FyvaX7yYE8DlhWa5WaZfAs4yOfZ90DvhSUn62bYu3pb+5V4rIVT0j/8w7eW
FguxLfrC7dTT+XaEyQHNN03o11Rx5FXB/+kNlbBMHw4cZ5MzovShBzvWyDayn3MjM++vxOvl8ZaY
pv5ok/qPqIfg2YkEMD5K49aMISaj+DJc2LDAkhpemZc7slKa20r/DzHKPsF1Ki9rQJM0wfEmd/bo
RmPlnTjaozPJ/Dnu4GYsxk9jkUWsBVEgIGVZhbWKzEctRI/giu6r1QWDRu4KyFqC3hrNsePRkzJS
siEeiWfSrhmkIgX1E2+Rg86i/E8KvSe8fxEuCSlBfSvo+ilwlGWh179MThsYnU/YSaVoH2FTFGyx
jdNh5822SU0HPNGMo4Ha0wFbWtVlSb9DUDb5bX9xc7vvMtv+va+mvXhyZsa56hyoMJabBPjYRDYn
hzOHOkQ3tB6koqk+ENMQc+s4JjmvJevL1Qwpup+Bk44Wki1FegJEU72KKYglKDlnXGQb1fHGkW41
QJ49QKodlVa9VzF7TVRNgOHhWikrjR9VYSX2+lh7ge71q0IgtJgBFjTNid7GPb+sQb8sMkMr6igO
OOzaXs0FRJjgRo97lPy1d9sckw2nHJ4klleqQQlKHCbUDTl6YHIs1p5U64NLcRDgkgZdgMpjLDXB
sZl8CVomEhtEH5SVCBnTqL1lv3/Rpko4K+NYgXFJW/pLO0/7Vj261qIoAsaXxgsaFccc/9cm1L6V
FRDObuAL+1KjN4AciXRf/ek35mg0zHGQAKJyip9d+ZwCWhsTPixUFBLigg7ZHL+2ZQYBeptqU2xa
IQB1RFnb+fkmtnQbB+S45QwoR0oE3YOJVtT3MlsdWnmIGFhWPrrlkVl7xMmHZKFgKWW/pSL2RVFZ
PjVeCKk2PdWezNNkFJ5gSkmtrlvLBz3T6Ax6oZAeCH8+7NyWu+nXTfLi1He7iFjl5yJGrwD3dIfS
M4/bjKoQFqGpeCYiBwQuaXqhV8auBt5iK4G/0iHqB8XB13YzcXE4bch4ecHmkHdfI28IAbgnT4Fd
87oAscANXH91mwO1LyiFnhi/1dpRhiELie1es/NSqYAI0PcKxJ1nnv8wPCG/NJcabM8LvEnTH9YT
KxlcmmQ0FkcIpQ2Vg5Lf/ERPY+2gV9uwFbSqA5IlvM5flS5gPJCUmLzotTu7yFkl/OmKP3pPp7Xt
9MHy+OVnJ9cyqWlWUct1C6VtnwnpaSbdcCsGsJyR09BVS0t1rLT3GIwzAqA7XHUksi6PbT+Ewgz7
2IazaRjQ4jfxIBJ3qPuV846k6uI1GrYm7MLPHZUM8WY/nxWgDnq2gPaNTq9O30hYI0FUCamNtGKj
el6fjJCMoOPAjrt/MZj+GmZOM/rsAfQLpbIfoMVXaAkqH75lkTecZTMVORP+sPMZNblonFrj+cro
+qMK8yIDtMft0cChbnL31MdlnfL6IBGyCqX1VxVhLah4KrzJBhA83AMq2BCDFwpUrBdFIRICfaIc
jF9VEHR+z6Vmwg6vLX5sVG59+JQYYqNgZYQr/bXE7mCmDLKHLj3yxvItoHik1yIDctsSCAwuwuTo
Eb5bS11fCptnWH71vRsf3r3aaVYewrK41i1cA18uPLpN/GQMNK8o0DuPFx9ERNnOW+vnTOktTMpu
JbDKeWrlqRdy6L5ihmAHvDZr2KQjDZKUCMfyJSgOExKvJiCQ7NxYR7toVDfhOD87jubt8nlfep4F
Og5tKFHxKaY1avzm5A7bHrUquZ0+hK0TsNcE/W/fCEtOxDpuA80rf4Fuv0umSlwLc0yXMpW19nJ1
zPCBlZgHYA3bd6wXiEvIpyEBUmhxLYa2BTtdPofmHDJ8GVB8PavICZOcAnBmCIKJ+adksmPp6pYC
x19TMtT4K19DBtLYIe9L3ZxyPhuUJ42lFnzSs/VDH+JMCN+uro/VneO3n+MG/W5sSb7WHR3bRLqc
DCyOIW9PpK+UCYG4LMzNbGh7Nrrso6Dv3d8hWRsC9qTxPNczIqN/Cqg1mWjyeiM+D/PR4/QS04Dq
BabebgJJV30Kc9Kn72vT/vRl2c8gVXLWyAvutyRs/O/J2EPKgM54JaFhYLF+c6c1scxcGg1TK+x5
U7G7fOA/GdGdPgKoKhxX5bLoqfUvdX7gNLX9kkFHosrYBdCb57x9Wda/p1M8ILIMLO+b1ALRQqYk
9HfaAT9SkdfKLGyd2GgHR8nSRfK5AHIM8sNIEG1OmU9FCd8BgvlivGazIcDQK++i309fPEP+SfUH
xiaoLNkEmo3hSWmkD8QCOSb8bgMyHq8pIWALriuwLffp7TxU/DRSywGebx8Xv9njOuZHQlAlo8ws
tlK+GmVlnffK6IvpeGi0/hMgpNYseFcVvKm3Crmsa7sYCVdFRC7irXvAZbNR9/DSRrjpDx5Xa12r
JJvtxwZl3quhJc9qqZLTAfPnvxkMvJEqBygCJn4lD6UlR4wNT2C+NYjhMEfOeGvLA7Il1elSe6gv
59jtkKOIsHzvkjgjJrQZabAgOZGXu+4ugm1j7RJHalf/HFtq6nhJBLCNgQApqz/JyxND8aA4yMp8
vK1g5UI0XB8P3g9ZUgs+JcRt5irDvBeyakZ0lZ0Ru6OhzBgoCJcmv/V+TeEHfNJUYXSYIjK+evke
W9h8cY8tu/t6o6t1TbysdwopejvgI2gDTBLYhSjL/n5N+bAJLb/0LFWxk/MPr/7rVGKaD6zxX81d
LYYUq40N/RiNXICBF+EwsWuftHR3GmecOLhYEpAjwQg3+cd/QsjMCYBQUWmBEKc9nJDObGyzuWoX
hy3OaiL+eOevY5aXFiGjOndBJ+JkJ4gXtIJirdebfuYNZT6/kCwIwktbK8jNhWTD6Hsg9nE5Mgdu
zYOuJdIbuL5ccZWWmrd76bRDt63vOr+oPFOO3zIXY9WQl310ThGOWp8nAyONtpwor12gMifiHP/S
Y0MvrsOyshHffUbiXikXgsqh9cLUa9R/D5gWQSSgcJoAYsCvcCTpDiusfNy3Kf71V6CZsv0xEMNZ
pIvWE+ItHOYRH8Vk5iKmajaIzewpcZlX67R7+2R11FKVKCSc37xxBeWjGtA76beoZ10SRHfKUvw0
X0MvaY8weXlT6m5IlzxqJWBDSP7a7pNtXFEJedzNtVb93kCHfxGcjHlMTS1aoIyLaLlrK55aNeXU
BRBSbz0Y6uAYEqL4RMhPtAFBjhJdt/PAw2d8OiHs1NjqrH5usIdtfhiWa/z3Zd3X8EFerO5KaJqM
Oe4g2cBlDk3NbK6LsAITR7AFAO8Wd//DXOs6cMdT3bniN38OfxPxYqlqA/SQzyoQwWZPODFXF0Eq
p3VHlpBINlyKApmabr4qZ5f6NBGm8joNJwqCxG0lk6QBuQ27qVkZTaqOrJP/5T3sStfeE5a9ktc2
TS/cG/l0mCyCMfyh/OCa3ACLq5gEOixQZeD9dIyAU605zuowKkwGK5K/wCMi/rWHRy+o1a5JtpU7
w+rz2AVIfBqpmGAhxyfmiO3OtqZHEGeBpAz5JTmjqsMT8PP6ERNZawQdGAfPOlClCTkLMzpm9Qt3
VKYyTprHq3Km+ZtJX+iXv5PWeLcFVuSZZdpeyd6EDWrIBCDh4rSBOgVCFbQsEgUUPVqzaISYxRFY
BU5a21W0HeQKv0+S0Cru34Z2RuKGIkSBlkOA6aYmCYcTpXe8doTWNKCI8971EpbJ8eJAHEJTFW2H
+L7xlY1RYs9XImZt0W1/nENKJ++CVEvTTZdrQcqI0JLJqCBioolqAjQvQuwGleKjLx9gFu46v/nz
2sjxhg6zkyS34BaaFpWho3AzyxWaU7fYVDewXDolS5GX8LKyGN8E/J8710rYQCosJk2dd2HTmzXB
nN5nSWOFX+E7ks9Vj/0sCiKm215KWe90RByS2VDxdllPSeaKKCVsNrhVam4ejZdIuvXvE4UsBx5r
Oe8sJ68BBVJM1fxjci+n8Sg6QP+zUvC92OTKoj6ft9gecNOSLZ+dYQ0uBSbnW0fzruO1K0gWuNkO
4ogZ5GMsv1DM2dGL3ESsExCJruShRbVGO6OBQQOOX8Md4nYBFseTY3GG4qBHxjGeYST5JDSqdPDc
nU4um2rwHZ8MRpORQ1h/FZUO1yVfkUZ1VsynMwB8I3zH1yNJ81sWt+PRkm46oNqPFDXKfKePM8j2
4pDRDUZVboHOMKmEypXfSO7p1y8jOQ7RM+Xmx188vblELa3rf9bQ5dU/LmYEq5ofWEQsSbkCygv/
9SCvlcaVvrJHHS8DpPToNMiQMeaZjb8UoZ3BGel4QeWZGAMZ0+pqhT2P/VcNR6xRsumiQA0VCZas
ngLbtR8AKEezJ+sb8CcBlH4F2m03neZY56JrVITLywvFiIPHR4C8YqerHzRK++mBLwrYdozHfHBx
wfr6HcxOSYqWaj4SQhOVvkrQ+XQqhdyD5y1Gmai2H3LtILUBFzDzUh/7QNNHFh8OR4zHg25nvj2W
97rlaWQ/y246VT+DlC0SCZ1UpIHRyxouK9ZuDYXcF0DvhytuKnNk6tdoUb4bXjjNfyswzx7TMq8t
B+KT+TvF4s7ln/NEGUaHoM8v2+G7M6J6aM6js6ZvIRinzMMxMcmRlULp0duwgXxfdtHpsDYzQ0YY
2RPqZd0yOYKmf43v6wag4Qgum2hC0GX4EmYPOtrqy6bScqT4lgt0HVKFzPwuoxU8H1o/TF9/u4sU
fbjkxAKWCcm9j2hyfeqm5Q7bp9mPhcfuM8d9GY+Xq+wpVMRpiDRxAqdcNs86ZVI85nfop5HJep41
nqTMtWdojRMUCMXssH72jl5fvhryBS/sMxx50Er8KB1dDuHVo7EV+Ow1EL6nqoTU+2FSKB82rbNE
lNfEq3yz+h6q0UzSRONTCcYaYNA2bYXgN3X1qsAlQApAauWq84kVN+Si5RmEjTApwNA62ox3RONx
JnwWhZxgFOwD4/LbFhlnuKuubjWRDT652LHGV1F8D0s1BSfK/lvxo6wRbJpEmv7IiOp37cX+IKmW
JZGZeaOKB37yFovf80mdTZYZn56/sPZfPCwigN44m0MeA9LGpt32F92+5SmHbRBJA6cyhLRBsXMr
6ZWNRWqP9nEwLoaw3Pg2LAiMa8AMbaYO7e2yFlDeHS492FYz3CeZ8T5x0OK4FnN7pP9WjNACnktU
OukLwn2j2WCqapt6jh0phq9AtnbYf0qKhciKfpjFNkITltroYif5Wl6zG3LEmgYVDhbJp3bxaKa6
qiFyTE8TLeeBXw0alJLDye66Ljd0MUeBPCyz09YoPlJXvc2f9lKL564n0MzY9nq6wgl5JT2IsLIH
LTJ2fL0ZH9KTedi26MSjsLpXvQ3b5lYKIDPxDonegWaxVI6wcvroO1be7nfur8lSTDcRbabgjMo4
/ihcbaNdDOUOkE+vN+RtyayefTNpQA/ycqpCQYioyLzZHn5pc4neVZHhy/y4qcIKGCuYz5FUil0g
Vvsvzbnhbcunt2+1dKuowPSX7psCconDplcJJUgV95diU7Y1UuDd4N8Ug7OzC0WLGDDCZcNpn2x6
3zYctlfRANDpmK291/ktDGR3Zy/82QAligNaOWJ/ZIamxmFNTba4ZERvvjdBri3hrgUL9efMrEoh
Jimc3nwtB/g3tOOksuJomjrdzeKoklnhhTtbc5Ycn+IO7h1Dmoe9+ohmPKWfZM1y8/bTPhvFI0JG
JsSu3zYACvChU2RNx0e/y2+vhSYUwOa/4y9DBk4z172r5nApSr7rWZ4abA44Yin+ep/p/YwdSbkL
O/ry9GQzZWBPGA4lAxAiCBInBnpE1RMNBKJ1PkcActMq2GwZCEdFP9KhlPEeAtmLrBmNNYCii0ND
d5DQxWDnRfaOA9ryir3gnFz8sLkJ54/hxO/b2hab07EIB+/U/vJvu3aBdHmPC7GVQeIif5ewV8iM
1Wd1FJLRS7iOJrrcSNaDGI208XOWVUXNROzsobBEX0tiuXLOmAmN4CSpf37EnQWW2aLcZLRTiFyw
BVViylocXykHacN8kONptoS6ffo/bVNtC2qj1D21s22QZ+Se4GlPd5g4idor9jBn05hDzhK8EZmC
y5NJVORfzz/vUf8gVbmP7AsU2p1ccPQnt/jWuVs1wBz/fsPO5ZpHDhzHbUi4hgCurpQHYiloWifa
uLD11oEpZbpGEx6CKugtkzs1P+rX8JDjREjSUjNLCdysPKw+OrAJvxQF8RFhb75vTIy26YUOTicx
4Vp60SKX7HspAR/WpdYauENw3334Bxftt1kvEzi09ZVjN7gZKlS4sWFLiPsOun90ZFSUlvrK+N1p
NJxZmxpRyeU1DT/zBVWGsGjm7nHtm85twDwbCE4e59X/5yp/240AxqDY1170WMTw40OKHTMjMUxv
ghT0D3r2u9CJ0TV+nQvbRY0CgJNzCspfugr+L9Eael4f7z3Lu+QB8ye+I5g17HTshUvXLcgRChLA
vAklTgkNajBkDnHGTqgg5K0mjS9q6jP+zF99hTs5SsL92rjAdnSVVXVJdMffAlaINlwL0JzgOqWv
+Nr4Qry21Vkz0Hxj9ri034nrKQoxIUQhPFn28t1RIK+XWAYQwzRa7lQNDKWbkmETHyIaOxxgAmHR
6YCVEfaRP6iJcBgy7Y8rRSgn2Wjas5iIJORHBa2LXFX/O9fcq2SCfhy+WKth+i72nCBQ6iTki8Yx
IL5jOC1rm+qGcoNghA5G4YVd2CNb4V3dPIMiXrmtdnMYj3Il9p0l91R8qttebYs5lcfXLP+alAU1
njmj+2DdSbivpU8MVjkvavnNUN+iC2eYpC8/eUds1MQnMV+mAu3gJBjhvB3irbc0kC31pN/6oH28
Btz/79rTSwfc09K/Lflctn7/MKB7kycBzf6LDdrC9qjaRIrnx+4ym/hapZvfD1KKaqn0cMNQVzys
7IiGCKPYsGpCzBzKTX5lZbsn5sCq5vxpUZXvhppp9ffzeAR90bNQG0eZ6O0oJ9WwOQdPhKznx/ce
4BCFnSbq7ZLYdlM0339MhHvgH6wRtr9jqlNlcsNSeaOkuzm/SojgjyJDOAWp4lkK39SEXYa7SDw3
cR5xZRiuaxLZ5Vjc94C8RUzUMz59F2lxjtUUOkhPrYoXWsTjhpLtyn1paZqh/BEV1JUDvM7wB+7i
wOo3yBAOW+6FhXGiJn+0HusJlIebBFX6+2Bsye5t8Sq1ICvcdKeNn/faHIZ1N/QxhHh/AGzH5PI0
sZH9yZiFor0qo6jheFtUurLMUcsY1JUpUuUzIHCr/eHA13/UCiNGiL586WO+fQFG97H4NTi6o25Y
qoXuMafZ354uC4WziTw/eNP2IYvbkAN2fCRhioUm0P+dCHn4TaI4iz1Mj5KRv6LE48VwZZ/eqwCX
iXLOVhPK8P/hbYf6j4kkKyefs0I8ErZvoPmVR6FF7NPJicDCm4KlAZ02lqH1W6nyTQ8mvbEy4ZAE
I0hG/SnXNdKIMb1kC0SVaEJLbleP8I1C6U8/djozl7lF0deVraWT4Z1uYSUwaaC7BMhvtFGW4y2V
65pECSbg/b+9Vcpt4NFvUW4BuywRgiVPybiel5iKTXxHCMJPsiZaRVGOFhydHmjudbC2gbdC9BP+
lvhEl5YXIEXRi8++8GkQEA6rinHcldOqp19BXl5o1KnI714wuh4aILICOmuTGHUBCCuZI1biXauI
EXwTU/jBnELW++GcI/uik4BzvkvrznAwvg3OLWBdbYK4IBt1UOgvRqeHGmZcyjzaXzODcSJ5BOyY
Lt9qpDL/2TVwgwxhPbp4FedoF7RNq9Oh6SCqHZQLrBm+v2rH+FdBowmg9krBhaKAmaekNrfVdld9
mFF9/mlsR9EXHa+JvZnO7+FnPyvpu+BYdy89DDYiq/5bY47+K8YxzlbajB061mtZkiMYQ0WfM1El
xMA1uPyOKSZ+x3EwyMCiEGuqsTQP1+Y8XEsB5ecRUmBD7+EAZqS0Yvu4LRJ660sa1KRhTY7nTInC
SXUO/HnmGTg4Bn1EL0e/rxW1hDPtNejghf/cx9v2aFmeCx1Ms4RbH4aKj8JouQ7Vz967iiJLA8Cl
sdHI73j06K2snhGsGwroMocMwNVrW875TByRTSXtoeWA5u9zd4/hpx65G8k9nlqJDQifub0Zy0Wd
5rpK9I4Alqwii71k4L2SH51dw4jGDlBlV2UBEeuvIN7zhvGBRgkEvcAIHZvkDeJwALFozBUiTKl4
2/vr9MkWgG+uZJqn88cgfCFFMDTaGbrupgjqW+kF1fZvk9krPpCoOKTa/k0rC/AhDsAw2irPk2MJ
fklab+JEK3pPrEC1jCklbGW+uodB1zts1bP+2e0wDxMdbMh+nPtaqgEN0R5RLewkHV1/dXYwGS/x
2CRu6gEBKxjg68aSlbhfxjCstykMIG0H5dNPaM4ln3Imc+peULpxZeGW0XEZHEhtVsYIVZVrz/CP
vz4BXLtjyU4uQIjDFav63kbwc0E1+rsQAYgMd5d/oGti0cfVEMUEbC+pkI0imJo5TLEJAzD0YEPN
DPTjNL8CjS4btbi2hij+0bjQIfuD28T3BlacpBE5b92yT/zTmqbUVOKXytk3Wv3AkhKO9kiPi9Md
2piPJ6cxDvQL6UCgfgFWZPTDVc2QPv4FlooPZSUMM2FedHEGeuQWUV/nzpS2tovIV7Cx0QAcgWa4
n/AUsKY8jLxVwIddPOE1VM8uMl4/A8GcIr6+8GcGbGNWLZBsk1g6RJ4JPo7oV0oxLLDiUMddCSRd
I/m3ChCDTZtiLlsBLHs1AAWsR/yErFZlMqWtRfOuNSpeIo0AQAeKkYNIIL7uYwMNcyqo/mmytVv3
PgVm4WiR2cW1Q4y+Odmj2XUhpfwJ0RPwKQZnjU18TvzXK0KApVvolxGfH/1IjED/WaSlalxifN17
D+f02xj7OM8CONvMUnaRGPTzWQAcmTfz9mY2x5xkhGp/ywBrTYbKi+gGmuiMucEkHCoZbQ4s55Yi
eq0yg3PhVCUatEjvdzfOJ41r2RJLW+WoH6g4kfsMAgnfOildtaAghq4nyRaNqsjAmAkv2/KleE0x
GfQRDwRb+7P5OwCxy9/tGaOMTItpEg9ai+vevABLFSL+3PJgpSVBxC0BI6i2pAXqkbfvhIXG8Ze/
DKrEhsEAMvjbV5EnXojx0+wu5d2KK4pO1bwbDAqcj1sx+c8LgxiFA6dcEQfv69kWM3HuGCq6vJts
kEUuDIvfxHSJx5uY954TojdJMXuZM7V7S39DWcis+z1IIHHgz2hHG5Zqq0gErHEYKfsCKHn6KHWr
L3pP7rRTRzciRdWxRb0ofRwwTuhnWns0U+OJMQzEkv7QNsWTEHJHNTiLP1faBYSwM+byTXaH+QbV
8EUWhUc3kKLk4TppOjHXcJqTRnJs42Z1vfHFsjOhHkR5fZd7Ch6qVyyCEqaeKX68jtK/0FIlNy3y
07tcGxPFxHihUczwrD6RY6D17vIrYvripJYmmH+7X1nXKzAbc3w+ADbMITJC8vB7MTSkcjfx2keN
vow/oWH+0IDYx0Ns1djsXTVOuKS8TztGiM4/E7g07ePKowveH5FJuSV2GGXvjKRgYR2WI7Q+CmjV
ZBD2QPdgp0xp2hUEBboZA7b4pWt8cNMvMNUyLJQuMjbTIfPZi3z3REaIGDOG3GyuJAiyFvKd6G6m
4CnXrbkAgfMdn6CkDkANBiqUy9unqHCIHIuDAYEVorIHQUrae0rUJlpppwHVsGz65ybXFwa29PBw
ajOD17QRUYBuXm8JtndwnTqosgmckB6HXPLNvfiYPFZnjO2yVum521B3//pMrBHLTinQb7ze6F9O
2cHi8HMwT7wySJWy8KSlFGSlodkCiRHzfFfaTWBTDFMxA2Ls9fVt5r7IKV3LHHTsQi3OLgjmJagS
LEA7YwxoLVnEg+hBLskx9i9cuFgTxsC0myAxU6xpR8mGhi080G0YVztzvaid/vPyrHTr0089A8pD
vXtnPOGzPf4VAnG8gkeZro69CqaAZXQtNa3b9zLJwpyDN6XtwJVEExEmYcLvBgiAg7eEhjicQshI
QiQtKGbJ4h/9nP4bK7BVvxhMOC3S44ZS7G4YvVFJ5xPfyY5IrmmDZVUFyRrj43yG1br973pF6uIM
xitCprrUubCsBYnsrE63dBhOa4rmSJhibnjKdyhcPhSNlpg12PJ8oWxa6cbFygNT6b1AUQnI1G+3
CKyEarjZ6O4FvLbibWO39UwrcnU6/8MQzqlOYpr19M9giijI/xGSmucZIgYJi+aygkRrVSAcFohL
ufIP/Nmf/rVULoyrlT4o9pO+Ydau5/pRRFsDujMxVqs7GioyFOapnWUPz7SlkEa10+prImC8hIU8
3zQo/bkNoSZQBJP5YxaPwW17XAI+gme6af8GKeGeZ8AIjObR6wiEdADLQP8Lz1kdg8dCxmyTYHvA
505vwSVhGOHP8o2SrKATespMEdISolNNauJsbbpUYRNRlLdymbMpv2Y+guoXvum95/FgANV9aKGX
fJfNXnVQAX5qI5T5sS/wRKPlodn8pFb2Xlp7Km6n/hJkPMUAfSrSW4DucxxQjTqjxz/xCrStPBd1
cL3Qqh/TDuUcDikt++Lh1mc99BW93bS7RONqte4VcU1LzD2+o8ik/G3bxDdzMSQLtN6XLuMhGXvA
gPiBk0yREw0ceyTW5WKwGO/vQvNMJd9atO5pV0xCsl4wHa5Z9zlLxDGui7kwvq9crYyhKcdo8Ooc
wvywfWPUu9AtTcWw6MJSgC55K+MUZOpXFEiQxoPaQyP3znUXKetIW7dscqI0y1nxtCDywLaQkPfc
QRjM5y2CCDqW7/O+6lIp4k0fojl+m+GTOVhNjxxQhrLfSu2at251cY32fGObAKM930e6U0Ekvh8t
6Y/uMrKEmFKIwlMgUzwz0wq1jH43QeL0Kzz2A911blMwpMpnnDbL6NQY+XzajmI1Of9v80o8R5jD
UB31b91fX8L+k1KGTAZfaQ3P1gjSnAbMFrc7AgzgHtqwi6qbQgN4Zb3bChmXK7FM0pyQSFxXvYEc
/T6vPFgVq05T3uthmdtSsIgzBS3oWE9FIlotd1xskNinX1LzVqAlNyuQ1FrF+Hxp3dm6ZWUa8xfM
RtU4q6axy1KJKaFr4JGn4bsZHoTg5DJWN74RUO4eP0dSlx3PjI+zrhz79fwVGrEr07Fm/YOo/45M
FUbMWWzCR5SUE4DGrD1SlCYnwo5IhScXOYMYLlSfUz7eJVEelgYFcDDMpXDKnc1k5ozDTLWJ/myC
hdV6DQOQZvY+ATxumwg/hbKCaZMJ6yc9EVZ22jPDHKctzfbw4A54lkWB30EpstYQFcjH2sodLoKj
O3G78cEvGg8yfvajPF6hMrFylKDNoLwrKGihHMeFq2RvwXTLD9XIPbQ76o44MNewSkEgCJswlaYc
ymrnUv+e2jyJ6wPPdCCji1U2WBFBkds/Q+1nFRk7E6BL6q/7wyO5sKpPMxHuY4qL9LVlNPINFPcc
+6MokwqKLzu45s+ZHrT5UGDY7BQ2hhDN7hgwF4DeB1/Rp8ujqQTeWTxr/Dvh1DYjIZ70VMlAe4yP
rsra34Y7r6aAOODggEfPYu6WactUrOF3dJwdS68zKZGszyKOsf1bvyvTbMnhOWK1OSU8QUrOOIkM
UcuU2diu+28SyoegBArycI5LZrhVTN0HTP4WLhk8hu7LiH1uRN/pJeqCIxq4/6SoguVECRL7DSgL
umBb7XZ/DhIc7AOlVGq0t/lpnvrOy70u/J+7KYpdlFpWsM63oDsyqTzd6pkYILbxoCt1BW19CtqC
urNccvtyVBmYA6vFHrx03tKTOvnmzZqu3LhpubJElQZ8ya558VeM3CLzKQiuYFbc3CKjcRoVDVJA
mEd2tXqbbt71bluZG/MzVDpnZaPrNoBBLYE3JzoD/EsD8NJwC6Ad1s6Bodnn+2WvlrRftgQVg/bS
7xX5GdfbRQQHv8W40keiD/VEUr3hBZmBiMkoQEqV363FSHHrY+Ypj1RsHTdCl5R6kbGZdwEdCWTw
xVQ3gckxajtwCM2iO9gs/QxI9Edp/UnOiPn0AQlGRS8bHRgf9fpUHBVjSOImgQZeVVM8p8ZmmBSA
H5qxR2AMSI4x+cYlSz0kx2TLk26SW19ADwmOGrjm5AeI/bVUIwcviw6SHQDxtpTnHISVnihhIqbD
+ESn1BVg/BD/pbHbgb/gH6m+g+koUOymn1BRykhYWBGu9h82b99vvYzRIiB4EqKUc37l/Cj+7Of/
vOCHZOIfPdpJlQl7DXoumFGH4dV+FQeKQVuaRKPtemy51L4HZUgkV8Svb5gA5dca4PZ0fmrW/I8z
teRZpG/E6a0gburN8GSBliE5K2+3FyiyY3OvBcJwxgGjhawliwjQ9KSTW3ns5Z9ojHGI6Od83VLA
urNU/grHa9Ar1IbdAyKcGWUlChZN/fuDNap1kzaeXLPAsJqTBjLISriM7CeJ9w4TSP2QfAgZFZaB
vXzVlCCnqa/AsAa3dFJQzOV35aZ3RkiEqtciS6dbI93KHPeodzkD0sl1wmDUSP6cC9wt5LQsgpMd
c5U1kR+uHfZeZvj1yP59vx3r/HGz+SMs1o+Q+Aj717MYKGKtpYzL8DsWe1sbllJLxB3jZ6cZjcqU
Tuj8f1BtC9nJbrc3/3hNL+sgtpQ7CmGzHz0XI9LhDlvIzG1UmQgAhHghnPXSfn1XLbcTy93R8k+6
AFaP5T0C+thiTG718SFHsNxZmBthh5lmF64iuMf6Jhx+hX78xWh2Qx1yc3a0R5w8GAoCovM2wle9
LpZK1KYqYZW9gFcuQg0iu41vJsdbByrMWC32OMwwTMmM/tVMuzRjUPRVkdINVW4rCVdjXfqnX6/P
7KiajpcfUtSaC2p/HNCm8DypSOnuka+ipSnCrNBrqZ5cl60X1iggBYrwT9rPW+bDWaLYEYJwURpX
Qj58jY69rVLZFcY5Ri+uOzLGXFTG23zJ4Q5MI0zOQWKVRck7qSVqWTZUrv8aUXQjYkQSKLSdLor1
qfG35uOuvut3snk7YNAwLOZZVY8UFJIhReM/KxxNEeQOm1HRVaX4yCfE7Nd5FVJt8IajnIFJSHTn
nRnyImasg6w0yVBklDYh0K2kETx19MyxmDAdm7xoF1jvz6mKisDrvyRtLHBoOxZlGdnervSqWDI0
EdWhq/jmLkt9qDBkoKX9DznRkdm4MHQ5Aa3Yev+LCf9owmkwdjJ+DGD5EzKuaovi6AJWn+nGZPyz
XQKMHJUMVSmhrwJeTcI4+Y4uJW0JzgMFCsTw9Mff+al7pU2bhZ7Wq9MQEF5rdNqVnp8Vm4+EaOqC
6Wx3AKBc2sqrUacgMiMCWUEvc5XQXn8TgLILuCKaTSsS6RA6v+mpXy5ugi9rN41dz48JIbw7Bpj2
9C6EWkG08xhuxZckaS08tkAoQYw4cSBxykNHzizbUirAQ0cTirf9G0bfouXhvhB4LALzWUolJ+D1
zMG78B6szz5pi+sY3+PVEr98uQ2EeOQnTTU0qEhefpJyJTWJuAmNy7XZ9yP2tfVpkntValNdA2/e
Y6pacKE5kKbVsPxTKPBqSSbib4HXwC3EEha52U2gEep3uYpQyNwEVFI9b22i8+K8B0qp6AdRFP9K
iOrwRGvuzAS/dv/UO+6ovoZ4USpFyHJ6Bfo3vErb1oxU8rZ8yXO2Ggx0KxVY4Sh6jT9hGyIJICwB
2F7PWVCIdd2FxORhH2CUzTcNAcK3RAPtHDh13f9vwSdML7Ija/pf6QlgU9Smy/I80GFheQcxLu3z
OUfMyANo3+THvSrNhvB2bcvpQvHfLpZViZVl7zkEZFIiHaZcGSv4q+QKhnFfp9L+2boxP1tRgbOr
4OdDf+l7yGa/e1KJAPu+W2OD9/LGxvFMzawio5v8D+sFab1E1Xy2u8pU/Mt6vwy/sAPuFRpIWn96
N1CzzAdCkYCZIXLS/K1k6UxzKTtdt4sbYsS1/OBdssJm7iaLfEs+GBiHks6B/meX5r4DNvRterxS
9ZHkLPl2mMM/rnOL7SfoVyvZOBrgeTu+tKI5uxqkbe3FYTjSdztsFidqJxW0py+/hmtTuTs6eayS
TBaAhBNS10loOavReOaC56M1Zv6lDlWwfS6CByGWRV75TyApfh8kLiPdKsnGZ9twg3s934ydWLfk
RBm5vJY8B3cwImCIEOaFFCUGUhJjfcqVTxtybOpPY7j5lB7zT5N5a/A7da/Hm7HWu3SKErd05zVv
YfasoyOzPY4csH9upWNVGUItWWlLnGEWvZA4qHEQ6wGf+8WyWj3Q2cWpKJV522bqjPfcpq6FbXaM
l5KIIZGdMd0VK+r0AyUuTUaXdpeGKkcu/SJygJgD9lniIvOsmXRfFXXH5WYAw7hZ8lGd0PJTz2Fp
ivF9hdpigVkZTQ5zW9kSajn6ESTn6EMGLT8tFuHBLcfcIVWrtpaSwvh1jwfZVawDD+6EaT2gyPxz
iSJBHJFNJNNmFon+pLBXULNHbFhlOOkyqaQsXl5g3YUYLP9gu8wzhcQ0xvyamfTvfWuFjOo8mJwZ
TYU3L221qlOlQCvwZk5wE4eMng8b+FdWvhUtV7Z9lMg2Qor9XYnXsKWZuR4h5NGyywoCJmNFTwF4
R5BKMHJTIEWM25t8pkKvBIhT4i9Ke3H9VvO+Bnvr8ASLqYY2G1ZARhKyaDtKYDDNMW56hKfiihgU
lQ2wBK4PTlYuRFQkRcnwWhc/OSdKeb7c/1f7jdUXIk71UJ+IE5Cah3ew5Koc6n3owaLNxIHz3q8j
8eMJpywuhD9H0stPARbIG8X0mNhdVQ6GAnkqpCpnIc17Y0ck/GShtYk6L7dtdcjBMtqE5wCr2RtR
A4EDZuuflRjTVgNYxFcZsQ2ebpyGqxOybOJmPtApe1QWdo2fSUZZ97vWwzhoBgr5rHkpRnsXCXUX
2UD7O26X66mOmuKS78qN2xyBG79UN3xdTNPGYwR7bhs0TRYKteWrRWuy1pM6IiaGWjxivLlsIp4S
Co4kBw8/8KS+jX3n6v1x5wlBF1FQKs7jq7xmoAOHkeW0bAC/Fzj8ZsvyuPj1+S9ZR5+npHoMiTp9
4EU1luqVVFyYbimiRD9vydsqTbJD6MK1pZXP20PxYX9044OYFgf7hJrnL0vfdl1So+lm5+aa2FK7
mk6cWiUIj7kP88liQSSggx+rJcLEZyeKftLltSoyIeci3LvXQCJ3iBgztZIJ6unr5SNHxYCLiOkp
RNCgbjjvd9GyR3AMeJd/qEG64EUahFW053nFCvWhT+9MdgHLqKvE9idiZuM5RYBbjawsch5j+iSy
93SNKyMH2EHW4eLyu9UhlHFGtqaQXpWU+clvZyFZjq4DtD4LkrJwbbXRF/INuVAnPLQOyg6/6wxX
VDJAuAZLqYl8RX7CZvgXFjCZHNo7qB8eYFxKN0SAwS9ADadX80/mJDVgm/ECRKPU653Pb/xEvmFp
lXt1Lp0OmnrLiDAPoPRH3d2CKhbN7eoEpy5TzCRGp2fRD84S9G5MnoJFoioGzvn9Yr+pGEOx54eT
o1E3yLx95CfA7DURtBtIQKfhsGDxfWnGOvhH9e1ELpRZ0z5jtrvo0pCDIL/ecEjTo5azEJWTKy4B
jzCdlJ1DMzquxYA6r0V8RyOnyPvA2NCdI1OGtly9CZZ6iut1/LYq8tFPj/LXJWTWZho45UaZKPMN
iIMpebUe9Nx8iqK3zrP1XvKnPDW9HvzHkwdUIZRPDWB/wuKJtNH33zWtRQHKUJBIfcv3HpihD3If
/wtpqG0WDpopo5i3/KXlLrJWlQA0fhSZGfIYe13Z7+i8Dv4Brdlp2CgncerLf9kI5EQqpiujO606
GKLPvQX6w6dfv3qUAk23c6iMwYVvTxOllOoMETP4G8Y7IwYcRBkITZD4HcPjWzvzrEHfFF7jTLRN
4zY7MuBxPnH9badtyJLalH3iyTOtybcwoQuQ/fcP+TUCQpKXd3gcenbV+FBCMjPxeYcRdILzis6y
S7gg5BH+UI2ANP8KkVYq9yWH/n2EeSzTbUi0FAyEVWduHC2+HhRL/m0ZX1TE9s0y5krVRSs9xjNW
wMfsmfgNuJifBP/steBljgupnuNt5A8CTeuIH87YcY1BEATaSMZXOzPtGE099wdouQYRosUd5nHe
379GV2wNujVGuWk3kxdS9NTpDFwRgI8YbW7VJo4msnevHkFOwzh9dBwgxGX2g4Mpb7mRGZT7FEBA
ovFcfxDXfxiSrByIVLzQ0iC3er/7ImS6/3kptkyfMnOoVoqYdDnRaaRjU8d7w0s66UufYs5/zDad
gzNP+hTniVLcyFi1gg/t+Qmeo2aaM7AI5KNngCuVWEQzDoar2f+kABSiAtmcn7DNJmahJZLjNrFE
VzQBn2Wbwarw1A0g3SFkbgxebtEFRaqqsnQpznf2fzg4mVu+WetjaCBIEyBKbDWEuyt7YLalWFmj
g6lKAPMLA2coXzU04Ex6xMoIySegvIJHmHYg36qOirTQ/SLpDRJVVaFv2AaScAV5ujOO4tLfhC7L
Qz/8kuN4wxL1in8REOanoyp7Jyn+5/tLbJGMmgQEwy0R51yARGiu3iH/Qz+Ety47aHRnErxWHeR0
JMIclhgrS6hvWMwZ2xLEJ7uYjgP2lf9wBg4SW/LOGM9fjn77uyAIvVH90RzZ8e2Gvd5hEclGYNVo
32l5x7c9cZTaIX8/ItA7QDZoP19CnjqGMXQA0wgkupWbyD7pk9OWbbqdlNLKgTPAbLg/JFzrCIa3
3qWxJW1jJ3FAtjnvkfoPaDYTboXw/Z8BUcYS6Ss45U1Xd4+LHzZ8zL/YXa/fCjwLu/vv08fl3sKl
cylr+WNa+aemvgGd4tZmn3L3F9AJyC7SEd7DlYcjrPRUZAfpl/jykkDL+lmmNYvuz9uKAqlGWLIE
UxUPirTKQ/Jnw0sdjuW1UKPYVHuF0z87om09jWe3N8Z1McxieAEQqWJEeer/pW1nnst6KffoP3V3
1piPcmKpTqTdk72pk5iXju2lVOJSF2vEvbdS7u71ovvdKMepBJERgoiZM95dnORzb7RyWI6/whV3
4wYa5ckCCMXJ5hsqGOy9t8WLakV3wK+5bxfnmMPwWNjGkyQraQyifHVaHBTNc/usk5Zw9XKa3PhC
s0A3yTY7GKUWN/BkNCwuGsxQ3g4q8q08NP8w3ivMhk4TY3CDvTBZmc0Ssc3wV2oY2w9h/CAeF58L
8fdUtjDml5iKk5p3OFrz5bx1BTKF+AR8j8drntw71vgsHmRKvkjvAxixg4fuM1rw9C45MiF5GDCu
++7BOijB2H57zqeI0k0aKor3N4aLqRHo2QLzUCQjioRg0wQCCaSzGJxYgM06A4PpOLQ894PjxUd4
Ux9KXu3Z/ZomvLM893XWBBptz2shnEoaIyWhkUXt1tXdqhh32UKeHxOrjnBzBExzbcg44z1DgMi9
Stn3ESwsxCcjEzgKBQJe6fonbzJOjnzGfEJdtMBWNlCtMUkDwPFK5/eq+FBM2/nCYSweNxATDsrN
8JCZYyv+/2A1oph+VXxcqnFlgTkzn/KHqChMDpO7fNSqpXQgMF1WK3j3O4I48H4m5BDbqNbmvQ5G
5VFpkXcY9zMxIBI24NBQDPfCp0L6hE3oVun2AE46fypQqeQjEu5Q7umcChgen/zdlk0w8WOs7tvI
PEYPPtb70GS7S0zQHErcUg6+qUEiM6vygvHikXRDcqsj6npondIO/tFeoXafw1s6hADPjZdr6cjl
9bqTKa3bb9uJb001YRPeOsmszJem/m5dbI4c8Wdu2mNX/AdVYfGQanG6v4TcwLj+Sd9SA/YSJoLZ
IGVQXGWBANQf3aX1BiT+KjQnElL31QM0SSiQUahRgHjjaSXW6xQUWDmihCex9Lx4Sw7qbvGpsrsi
3IGaAJjds7beg7UZj+22Rh7qzRKa7h4wMBzww41s3kI0XA5x8424wozFh2TjMuekVKxH3KWC5nEx
6UzmopJd+P1qHVitPkh1iobs5ZlBnsQRX7b49fcHiztpu7qBm7nA0DGC/zLnfeISKq+u6/zqH2ol
sXEY1yHGsi1jCmpacTakb3Iv0JdAiTTfw4rc9UOZflxAHGROBnCJT2xOrqo72yceOBhr02TNyksj
9n+MuV9MGX7R0TuVPKtdA8D6YDohPVda8cxML/3wg7KjGwiryl5o6YafFilhYMV12+J5V8Co3siU
UobEZNhRx7AHWPfgridvruC/LJwZwus07S+f9WY8cj5UG3FfH3nXIdFTSEmPPmBdMIwS3WfQEWXf
SKIsor6RZkJ0lc2MrH2Ac/ZjBDxe4q0y9vlSNSmrv7d3ePHYJ7JZjd7Wb8v+NF3cM0cWrN8ujeU2
iQ/5S0J+yOkKh8bN7WUGRUvyhgczjiYdmxi8KalQzR5r20oXcGyhxKASiBfXaZkiWcgIsFUZh/Z8
bzRGcQQtqjC36wjuMoDV+nh2jl64Y29jjTcHaWdmsnlVO7/gEq7eRNdQTfz2RXDTrjneElOc8bcJ
6boW6sSpppdHkitJ1SqdCZipdv9s6fCbYj2B5AcXoc9MiZmbklqqvT2ojtDvxb8W0C0P/ZbB5ErN
tVtS7/wcTWMT0xpc0PnRwLqHUo3Cmxrpl094dLTycUOki6Y2zPYMXYEoIXlJRcyzQCuUOhzG2Hwf
1vGGvLHBhnC8L/XghOz9NHo+mY3mfAFaXaeFMDVBi+CRjnTZpBtjpIn4QRcKHct2SK1Zs8Ij1MlT
pwa/3VjcY0PAy3Z1kSFOHON4ZVcV87ViBqu4+dWrXqG/mBNqa9jXqRSk8iHIo2zyMGW2z3ZvN837
QHtGs90UdrJ2zX56pmgeWWn5neitr8JAnxzLtHPM+eL2z1J5s9HnTsBckbjkL9hD4wAuDzS2oXOz
Lx2z1TKFNc68mpeHMV5HbLglLDa7uwIjPS3WotAeqfLtS1uRRiDFaXIzJbrsF1s8QBIUG/rtGnlu
fVGLLKBkwLS99eClA9jlstk9I2/jnhzPG3gHP+nuOfrHe1+GEPZQZbXzUPMpv9DtIQGvguU2KxRi
TpfFrlV0fRJWLHFc6CVTVQAujUP2yXSyafJg+XyJGIFSBogsFSVfgPTh4mXNuJm8R5Q/QHew4rUI
HeZjCpRixkUfdj5fDgbmrjwSZ96l3hQI9zOymLV1pB1KTBWzInt69kOfvJY1wbfL/AiyfZWu9hwk
IlAPhQXVxuTaF6mwwzIi5bSrLK9dibbQ3ZrPJT4jgUs41YlLlnojdSLQomIxsPs1ULiuMPBPWfTS
T4y6OJQOj5E+gUO+yiW9Cxz82yAXCFxkfM4r/dhLmV/XqWCJKtCK+Ksgy1nbHLvpSbw6v/ZosBPp
0aOwjLyguL9eRF6bDsY0RcUyyrw9IlWOvhFd6RbOy/B08XweGJFG4KA0jWd0q0xP5Ncems5Ijoar
DMHGlmKecvMMiZvcsQwCWN80FQSKidPkdLpt8MB/i0sZbLlHd2J8yXapfPUizf6KI8CuxnVqmPCx
7sfZmzk3eDTXp4e1jQd9bqFdbxziduN4iSQ4NnmTrfsYjQJSPmUOSquT1znJ5jsQ65Rwumn1Njqg
kpef30eu/qt3bwSYpt4mbYeZvYdgABItm3Zu1+LsZMpuXhbDN45Ib+68Nrhst8YoGJLRaCvRYlkY
VbfwuMfhBXLAXQLCbY1c8XIZG4CD6rnhiBJxZtSpVIVmZR4QWHCmsURsiXZDpvQk0/Y33l66q4dY
JsACxqLzNHI7BwrZ+JuaVXmQF+dYsGzmMtGGZExQj7qho5uUVkjq8ibhicSSqW9HpTOACj4Zxnce
9OtEtY18Q0otcdF2f2cNRQW0WzUJWaEuErJWH8ocdXePkpyq8BqvfYxsWZSe4OaDYJmsOSPUSOtF
Yvzh3mqTiy7Iz4RCD1exZZR7+6SO3F14T7Ab+uVDQgRUe6j11vTsC/aP2Khzjd2ruC2CiecUDFhM
Rzt3UGcivIoe/aAGAef1hNFVfFxAPmuhGmuZ30C++6nhJwXX6TyOkIpGwOS5Dy3o6IUWGLdHPY5G
owTMENPG+L3aUJttGWgJ+YnuVt+wmRnsjJ8DXBJJG+iPYcg9ONqobUE3H+I27HIwkJavW1xNA8Ef
aGOlMB87Uab6XvnumVN+r8tKJPdt0cULLLlijUQLGGZTuiS0mGppcVkigVTOVAwI3zXCkXQ95mlj
2FjylP7JdyotYTYL2ZaKcuuvHeduf7rg2yApcc+HaOT3dM3XhAJuen55RSj7+5NaQLWXXaDoyE4T
dBXRxb4hE+RFbtg9kHGfEPWhDaKDDZ9kN8vAZM+fb413UoXTn1m6Zai0UzwHbWd00i+bVL8jsNbN
SpSkrSI7JcNMGvnnHMs3pYK5M3n8l8DjPD5/yn76j9exV5r979FBEKGRjN3+DWfLgvHaz+5zqRtB
y7jCaAbxJ4az38czBA1iT/Wy7S75OH5Jgs0ayzMxHEbvYGWGuCEqCR8Zt5eWz007SZPyhkwvpAJg
OHdW/JAUHLm9za3veFRg90QcX2vid63mWNz05iJul4kxZO4+gO4kf+fNWFxK1igvKIVgPSmPiXNP
Ik3ZRj4Dbs5k0d4sOIUuCd4k5haPvxTjbfCS0fSlU5ZaSq4vsD1az+ysVBS04+kVWMAkicEvOQ0P
FCyra7H7mUtRh20VW9K3VFawKbBnkbwY6zpBNRVZORaStPxzC4Nq5dbkjRIgfHbBY09E72TbwyJR
hoSlgPD+O/VCPZWZoV4I5SX6Scc7GKTZ2mF5TTQs//2JyBKkhj+w6ke6tqlwnAEOqSmspUb65lUZ
y/ms1t8LVbRmZdGhiU7XB+70K492OWcaQ3sb/mnV9EV1vGd85G+VS94tF+Pb2eyPIznPqNxZedP6
/lSTHfw+aYHlT4/gi2oCVbyCxevyr5TdPYE69LHdWu1jwE3Xq8rZm4JJ71+NZRD33hqfjhwW/sdJ
FkOPKhx61Gfj7Cp0iPP2Bue/NEveZkEe+29huhjWAqHQob7cx/zzWyx1aIL5DuVCfcjxL0P5YRM7
4U2pAqpDjyibU+xhsVnsNhQwxRZTDHLyDRnclat1FrmgbWVE40C9QxVk4BMSEO0Lnd8GQeLtvYoQ
WLjczXZQGP+s5k3lgLCl/D2NgUf5oSTeNLd8x/kZtcgkN4WkqeBZDjnTftNUevPFgEPv3/hUOMZx
GbwmRT1lmldYlAbwOI+pd+JlPv9i4BZquy637QbeseXuSdH5xOWKsA9EsuoeXNzEVami3wvn/TcB
encWOVqTi8ZdOCQoDeb1SE9m7oF+I17Qwq8SbQBnz41uvx0lekPXd+x3j681bferkGgBSFU+LrWy
7wPn+4zNIgXvv/tkQE9ud414SfHSjaXBvrFTnmHbhSx8a6INMULc6kT9cBLp/xu9R57pG1pbz4Le
7UaJMYdp3tRw5b4T7cA9EnkZfBDCIBJoEGPZkCwmAZAtZW6rUMHTxRNl1icM0tQfYPIg/5xeQS1F
1O7QDPJhra0wiI6IscBBsOwf8tCgyCwq4TXbxJNjU3GHYctsdYmWc9LTBpK2oLvny3iaG3UQEVD3
JGAGFmg2qOQzHH6Sb+7XRFnQdCP3qcsaAfwuwHhOgcoS/cGZVjuIpwT2LKz6DnJwvcJZfhfBjfYr
hIAiyOPBFwO7tkeI8ITna0e4Ahs3cI8jtYLFE6ZB2JiFB6mFTv2lcf/hglZlW3H/aCYdQtmpfNTR
0QaUK3L7D7/7nTg7+Gw3y3oOx8i/LfDD2U1ZVkLnF4F+ZaOdX/2l2h6GW/WH3vyn4iMFOuaUwY2p
yvr76IWyQiHuJuiicknJUDSP58tcbpC5OS82pm7eRosi0bPPhMjD1dPzZNp3C3zDb7cP6bgUeZx3
Y5ef6sXz1q/MNejWN4Zb3kri/HrxJkZFkSJ/brFuDPW32qHPww4y18/Fbq3XoxoGkk6NeR1DisoA
iHsGiMN2/mnVj0ynOFOCZHoeOBbYu0rEWCs4U8rg/QjILlLOTGbD0T1XBBEUjlfOYLeWbZk9LxXo
cnE63mOOklclyPZBilJAGfdH8Jmx9zLmFRRVtnMZCJnW3V3+gWyeME1G0wxhzf3RDXAmraPuoDjC
u3gNqPG2iW+6BdoEbo0Q7BvDcmXbiFCZOi/U3mZlwNHi2So5lO600+IvXSfqzvVzKHYoI+7Of29P
1GmzZG6zLXpp0ZrM9zqIbZz00+Mlx3SuWcmoiIBdSwwVsWXkk1sAYC344r5d2v7NR3VkBIzYeWjc
WlGUQShuI3JJ34TVXKXOIKHRwcwBFnCfoafXEEuyS7i/DdMP8EVhbuxEKEO/ROP6olQmHX4seeg4
iIt7W8AcltiTXg9Z9s/QYj4yJF72UVrkqw3GQk58LvtaeEHNy+DO3lBmnHJq3x0imh0mdQUB7wn4
Co95EMZykhoMXxFY3Ak3RqV1WUnE4ZHGF3/cZ4SL7Y8MGxlPs0rQu3FLRKTZiLzjCv1JTfMNQxgV
rF9JyiCdEuGDibGu5cGQI7ruChsfkEXchr/LHwitVviWOquCGkkvoTufDO3aQXgVadoQpvrZs6Vp
W4aeS5x0a9PouL3D+eRcmTs1Mjr5Xp5ELsKYij67l5p7Erqvp5+lOMasjwRMiGL9kqnB2Z6qirT+
adIrjMJlOSD5BesVRA7XFqnzL80p+VsPd50ay5yMl9i7EV7p4wdne1ri0lA4EQ7NP5YWqzs2jaNa
g8stCgX++Zs2UZSDkopP3d4BOGa2LGhTt2DGXr2FsfQAXDAYALc1i5qmFYFufxKExxPOtQ5IjYEB
W0+QZp7GcTz4JdhWy/OCvafDaP93b7Ve+xQX/H6IiRsA04T0F9d50HS1ntIk7RDC021P9aGRE7TS
5sSPUL9r4gVgaYN78DhwprogDcVgtdAEeXLTjd3SihjrE0gTDp19gc8YuW33cEboZPW7hNlNZQ1O
tmLQmw6t0oiMMifiYm6EA8+KfiquZdJkHU4e/qSAg2NkAsMuzjdzjLkg0qS1xD6dT1euX0OrQSUr
Gm7m3wqf3QRcTb6Wjiy1SvmsdL56gYYcIL5o713DjPu6z1t0J4R/RYr0YxRGJK+850Rvvg8wdfum
R8rkQz1cYVxyanlYyEy99Tf5t9uLon/f2bMhPG1miXy7MIJU9AsqPoOHPqEUW7GTHfaJ9DVVwpKw
04u0l1p9FpUKUcLB3MEWsghiLMFf2PwJvFtl/URNkH3smcGNyX1QVn/eaBNJ7Wm47Dj45bmHMLRP
firRWG2xF38ztxayFEvrn/88CTJBFtCozLTsgPnij5C/9AG+FFjr6U8Be4lwm0e45alcmL9w2Y3B
B1WtGVqSfqJELiIUT4aA/NPKOQgfLmpB9tUUSTQFICTeTaV1uvNFBkZrpW797L6l0Y07VbNMQP/p
V552JrVRvTkLF2o7zKsipZq63WAQ8j2BbV+uSAt/uMKGMbJ6j5n+BcGZmyV9ay5EUeucL5poago3
UepC5hfBuHoIMWmURtKJ7AbB+5ycSUg3WL3GCWT6ixd6VX/1zczeMbs8ypX4tAcqcj1CG80dEUGe
H6Px9V3I5s1Y3PJfZvus0iD5EtRE4HYK00stlJNhmDWHYhwGwUk1KZMRzzTcFpi+KNZBeMrjZaJi
0RXpnwe5CTsBN2FC7+YU/qxgxUhXq0fd4e/weHCQptzQm1LElb+UK3DtBYgkq940UpqbEjSKVJJh
kgnLkB4JqHl1sPZDIRyJ/9OVOuvLPRR0Baz5kJpE90xYypFLg8s0OCkKrFqFAT09uUI204Ai0sMB
yRZHxHn7RL3K00RBagDdwBqgeQgkzQt7nl5EUK7bP7IToh9yERbOrpGmmfKE0JE9QE2hYpmWiA09
eWUYPXaDvOxVGp6eCaH/22ObjzQ+QmUUe5b4hlN2A9PCoNkjxb9rzzHsbes/NY/4H24DOr/Rg0CQ
hbfYmwsqMij4yOMTwI79R2tQ+pLg1bQm/rPEVedf/A++ihXG1CvpZCstkqiIoyqgE1950LWj1nyw
v4lr+5IQy92okT2i1065RWLiFsWMHS/n3D1xzA2crfYrfRgn28bqiNIUs0tjv9lcclAxkJSBkyh3
PR9Df56EpEuxVwj7sPLoeT2yUTQXN/o/WSOrKTrhSpZaEJTAo1tvdeTRbCFgzzUy66s6E49Lo7dv
5Mzbu93EU2o28wJsFYb8smMtyS+LiO9YmforeTd5gmw0xV2nz+4LJbMpAuIHwNdVJ411yZsIy5+3
Sot3Xo0qF5eBFQI4UQr7IybVBvVwi5FciM3ZHCctNtSNK1u5v3gHrbiIB5xTo60cCYZitSP95krP
pMYsFeuJQLx4JQVSfzKfja8TFF0yXcNkIHrACRW/fExSytsUkqihMtIUjFBx5ECzWX64QTnLKQcZ
yrT00kPMoxPoGAwKGyfdH5hbf9LsdCjAbQq18nQf8VNxfjOUoJIVnmxXYGPMHCYAqjZOguphSN6/
0yBTh7G4MCcIDTcG1Z0caquwlAcI07VIIdr0vcFMaR1GdA0TsK+an6HeM2Ws+x1wNMGwMTDjAEBH
VxbX/Z6udDbsPhoecFWAklw8r1/BcFSCVlVhaOcV7A1eq56w/KFhTCUWUwlL2u5SSfRmxnT/yPzV
IzsqKEFbku00et+VF/VabSzwyk5DvSAycQJ+xSdk4AoZ+Il945qsFGr5S20rdSvZ504aARnFdjfq
dfCJgf/2+tGG8l1JJVd+yqAYgigEU0D1SQ8JvmHXwrcC2jAjC5uiIvdp3pKigA0i1B9UU3vHx56f
7w4BsolgImXJjjDPLO3kLFrJIIfmxQ7Et7Omd8BY34pZku4+uh3fLkIT4StqeIMgpdY6Az8YFv2P
KY7AHYoc88/F6l1FFJragrnyQGYADvay+YgCqxBlVHCeLUzCQILq5hePBHGcIsflNhNZMbqM0SgM
VSrKjPk+JXZjSFgxYBjwpWau6cAiuI7Q0LuCrnLXKUwtwDyiTQ2636uDAmOy/PVn+Wjhuy9kH+Tt
LZBiuNlF/zzyu94pWRiMdtnFW8txErL69+6RP8NZCI9E3Gfj5GoyjwOg5ccGqGpEXzhNOpnqIOBh
eOsP0cQ7oBhOYybQPQ3GzcoRzfwLpJrkbQ/SrLnFX6Xz3145jDCdZrfLA+zZGyIIcZw/T/SBUz5x
1RHqgqBMJoFqszTiUVLilTvFq9h+26xfpgtU4dwRzThCQdt2Q1fniEmHe/btd9PaO/2Tg5oxx6xu
sBZkKWPzr/UBuuMu3Dn5YHlmwsZ/zbDun6eTyHwre6sxMSc780N6SU4yOFNK9z5k4JLLnnbWlJwJ
xCYyxWvnz3j5V8c/CIWYcePpWuw0ur+0n0WL7/4OQMT2qea3eBVb7nVRCHuLtzdv83oOvLdJ1Ssj
GhOTeFjgc4J6BI8h0Y9eFmRJuN7POl2OP2igunC2soI4upANSSCd+wuUU/KXJcS0iMt+GYZtDU5W
48h0mAzKMjosIeCqlRkBhkuFrQkyWCtw0Y96xgMokXkyT7Yl9pjFBR6wY6zCS5nug1D/tq/bFEYN
3ABPRL9Mm/q/IGlE9EF1wSlr9nEm7fU+qSgFC9LFyLKB4XbZyA26DLVxpy/58DCpA7rfzGWxC2hz
BAq6jShnGSPE1rnMDS1n3aHTAZj8sjjAnUjnAuAFMqxRZXIAcAHS/juBNx/Q6xiayBMHpNAEehxk
pKv1DDWG1BDEidl40kE1JVUTJFwjuRAHU+1HURsaAM63T9YTp0BrK37ELF+YkPmKHCpsZ4sCzNcU
FmJSJyTaYfgjczQub3UOfuvMtflzsYCgfFgYsZ/vdj/Vxa+UtrxAQhBYk88+YbE0aCyNWqqLMUgZ
gl0/mgMi9EHCo63ux8bokzIm8nq7RfKERP1u/FmGF3Mk+3wKi6h6MfB43YJ0MaOTqYOCVibwtngP
yHihCRGlTtNvwY5Fp4oeTuvYih5D5/7qm+LupRqJg9UBCxvVdBduMBsWivUT1EHsQJs833OW1920
snUQT9Gxvy/d5IMVBgmiV+SEWol2Eu1P9QrNPvgt2E3C7JsQoxuZGMD7mlBNvBqehx14/n5Az/7D
pjL41P5lbtDzr6WirxF3rvyWxI9xgyWtudiNSXLpcZx3zD34vrrdITn/DlLCsVZ9QDSBW+mR3VxQ
03/Bt42a/J7TLg5Cv3u0JwtP9au6kdRexJYvco6XjWtti/rqQgHBApwN73gUcVP2x7VDmyGNDniN
vUxWpPuxgbXxNdf4UqWh2z3ubDj762a8bXi4/v14tJxu+dteruY+erytteIq52VKgjBrFn/qw4Ic
tFZI5JXSuXG1EkY23OD/RvTuxJi/4usLVzd9dcF7ymN7gXyCD+ktyBWVAzNGItMorRnJEmWA7i96
YgP5+4BJ8gMLRPABo5uluv4BszXcdw+x01w3N8s7NfJrrvXLrrQrJ3IcHacI4ziALtl96Tk9zJnz
5ILpBFmzDABUAgfgDa1V/WgTpn9wLAUW7JuXTKmgHYXw/346fF9T5TzWW3/HwYzRDgDy6hv9azXa
Xl2aEoMA8eT6zpYx5SrCPw6cKDKf+CSToCqie8ZHJ3HipVWkoQoHYceknyPSjnqMVBtFVjIK7ZGr
po9Ra6nyFMCXuKESim0A9IN4S7WTzQ1T7dxM9Ab7DWyn+N/6KHMBiWSFcXYjFjW5rMgYmTYAbtnA
TZF1/hwm0rTYAxTDI/+rnl6H8A1kLzGgvaXZSMAT1xO7GIgbJS2HQ+1RDSe0nUWrVGbtUyq0mW0p
bDjHNBG9kEUHKM8zwgj+ONwwgZ4IoFVunk2WU1kwsK0X5sfh7YO0Z5CxT9P1e66IZ6XUqKsZVxcy
iAd0JazQxM88pc6P0POQ/PXvpMBK/YUhbxMtKJ8oWDw8xctUBsAO2RYNi/qffmaGPIGi92J6HBmE
Sgy1WL4gfyQLLIUyjfxuL0pqqrjZ0c2zmYgLWFhfcC+n+yPyex5N23btYdHAUwE19uwjlrSt03kE
MwR6z3B5fRmtpXq3Kb9XverNLzoybCLwp+3/xPptlw9SNzQ/RH4+x3Hi9l4oaEQejOaW91FWmKmy
qmfgsmV8QTklPbSjVMaO7jdie2n2j2P1nU4K8okOCl7tPFm5bLbajEW2g+u/HEXfQKhQNZXizxtI
hWZzo+bCO5hCaH59RybitO8bAn+7cEw9ePaw/saxkUaSNYzL/TyJua4/8fRW4+gkmN1tpaxSHbYV
4XBSzxaCcZjTEo6zb0ID9mx0rnY8EC9K3tmU3wkhVVW1iRE6wcLgrFlAlq3CoUd1Iey9yx8DJsHZ
aw5pQJxX97GQp85m+X1b9c46lSjg+q/vgCbxuNw0i+AF584xZiJXnKKbRHdBRl8mLXy/vGlbYWza
eet+1csbNoSQfq6KfEn50r9CgRjUCqENnEcKNdmPLeoNeKIWhUtkeqpi8Q8xhj5tnfSpMj6KbHWy
45+WqjrCEcEKWa/I+mudvV1eYIje7zwmpdyEa/qcALEYpPr/52PPOJU3dWz6nmdLGx8Kc8n08Aza
mH8+aj2ToS1GVpuuT2cRva0wxYS7gCUFY2/vvEglO9nNgostsDoCQLeT2Sbj+F8ucNTRlUsxpcsU
O00i6+sq9ehQDOJ8Cy+NHPXlwXDw4etFgaHiznWzRyINq0UPQuveN66bajHdIDJpqgB/E6sL0kLr
1h0u9Qua1RYqlcN2L3AibZiYvYXa88H6u4VpwVTwy1t446LK5vxVdDq2WnB3bgq6N+quSWtdcapu
7skse6qudiYVsmIZ4AxYZJbjr3wGiPsNOIDJfocUqKZ1isV7W/d58oS7Lu9XQgk1ZTgTYbsHgDU2
XnlrjVSkwu3Flhe7SRCvOmFJWRiNBq4NRkF6V2WFLxyAH/tHkatZ81pwxu45JDCXVxE4wM0sF1pG
Xy2QNu/NQNsed3ac3GWMsqStpdNC/GOw7r32qNq+iSBWlM5gfilRqhQ50+boPXasAdvzvi8L5Yzr
lI1NSLpkIE49v9eU3WmnN0mB+7jlKFN+uwShGm763GG9fR2TLjOeRYGfdTFYvqunQXwysu2Oq0sw
GHQbcnL4PVkaMTb+/sXl+JZuD0DsArrhdu/i/XFZSAeB4Lw7p4xJAbpStiq1SS97Y85OzEVO7qsW
I5rho0s61T/PnwywZZyqrCRjdYoIqgAc9hv5TOV/0vWuuMooPlskjR0bOuuYQKdXLBqlt3UcaXjo
mljPzuXeXL4Ocf5rPsHfkRDHJzwF+U9DNMH0k97/D5sw0EFKi5jiDzj4MMlGAbDzAQsHZxX3kwku
tAHH70z62f08N7lulzvsE1rYzU1RjmW9b1doFfN0MRPG/ynljtNVy/uCYEfRB2/9KCjMCXki9nAv
ygPhe4DojnAwecQwPQ0ZPL3x7AJjcU8i5HDlvbDT2gb14+K/84Tc/SHnKRMQNwngnSAwNsu1okJC
RRUcLHba0JnfmT5o1XpOC+frXosCy5FqwLvOQOAASNDkA44Tdj8cMWdET3cqve8uYzBUe//bKCz+
wDjW1TNfa1k2rOr3W5WPcLjQXa9F6Cnu3egC9+qcohb/6FspclPPkVxjbQlLsWnKwFc5bd1YYrKS
VtjO6gC0/b8bE67lTEj0r5QyuugwCZZl2rwtbsmWNFmZkOJqKkAqYwTMAh65ZGXaz6dFlZmgTAhK
LCmFzt1Di2B0KnKW6hjP7n0EIZBIVe+fgOjOUOtyNCSbXyLq7AHurutGIPUyZQtPcUhKtSBWVF/g
9uGUqLqDIj5r1OoBoctDqJ4FyGVcivMvF5dHeyYRDZeno9DOw5pmujcQokR9g2ndV8a2zbmOvKkd
vbKg8n62lIuLanSwLmS6V0Ow3Z46JmlWd4ZB9XQny4TyoOakAmnW6s/uFPjUvGh9c8dI+yuKTY+V
WfCEHU7velhBDSvui5QWtGmVHqopsw+piG3PwMpMjkIeDbmINK28yCVYYtSjVZmCZisrLRb6PHgU
ZMtPUy/J0nUoZq5IulLrS7Vl7lml6hcRMYahOKzTg2gvtAjdV0AvNNEVcDQczrzjCSqlw20s5wNo
oOEIeo8ygFi+fYBo1vlFa1iOVLAO+xx/033rv9xeUiVbk0mHlZPXOMxZKm6CeuXl+NLZAqFlI7kt
2ULSIG37WBPIYKRwNndHUDkI0Og687qqMbj7UOAE6wtq0VMPdj4u/rva1rzcLVPqN4ZzA02e7+h+
QlVknwy4yqy32n9ho9cgQQuDz72Kod2Nj+e5rD/KkoSz+WVNthBLiSiHwAmCvPISTeFzTo2YgiLu
7uBVtg8ozakwFV4sjxI63RrjCbKN+XouCYKgQiTgsz+Hc6lSAN1b573cAlqOYT5IUuYS2Yp/LHKF
2c3jrxJRo9jidO7eyU686IKTMcrwiQivjxhBA08TRmWD0ZQG7qA0NACkxIhe0T3Nb+C3Godgwhgq
/ckHP0e+dshvZ3wEZ5eZ1sEvCZ9l7jtiYSKwaMKqSo6nfMfE/m5Yp6xD18M0eniLsj6FSgkBkH4n
MVyGmcC/xIDzp9GY1WGzPfjfZ8BryUW3IhCus5tT6bziaRoy7Pc5r4uw0uQgBMbI84Z/LDQfYhi+
1Q+FV/nZhSFQWOTTfMBccUKHDtz6hdNViKY7rWY5YEUVfCzwxskhntBoPew6NfLGLMQN+IJnhN+/
1VmqL0FBdtRv2PsZOLY5pvzbSq1DaPOIvcCKn+IVDbLqBE41F7jwU7lQK7Lz1sSb/8+TsxVKunnH
4Tpy96qH+5kClZWv4ifMWCsyMmbxm5HfnvRQMHq+5kuNNHDAqelHAaSswRlNPykDOLxOIr0zf1aS
JhvibN61hZKeGyoIHUdfVeI7SwBKAfcKm9liFYZStWouh7NZjhIJjjcvm6uluCK4Wb2iV7ILETsd
8tk+ECtLdjdrnyL5E5JbQwv3YCifI60pgvJ4MpdnrJDTm0WxFaqWiYWfW6jYkGeT5mC6xBYfKs1A
NjHbFao4vh63q7KaCnsOp+V9mdNocjrIOKoCw0XVt3rwmotzWjG6h4eaZi2EAJNd91/i4jgjcWXl
CuoRd6gYNcdYa2WADeCBr8GrLQcSLzPhio8fukXPDbrnTb3CyyE2ROrJ1Q1e8z9etntOX0mbLD22
1oDtLJ1sAK05z8fHKe6qsdZtBa2ZA04LldrjONUI1XLyxmPfDVpHqK4qUV1LxfgBkIzD6dMQTt4f
YOEH7wxPdEON4ZjrTXWnOTuKUd8Oori+tnrp9/gtyX5q/g55MkmsnDLIWiiHrQx7TuiTphCoXrRK
EQj6ljXJR8E9xykDfNTVLu2GnwhIIjVyxyWYZn8ha/Gt/poZjgO3G2CsIsZ+Lo881SnryeGEn8mp
yV8p4acwn9H6gYlHnehnneCx3llR9V8u8NTzp6kVYvN2HjgCG85IpmYtf+Otf1LXZhPco3tkSUEQ
wMHir2ftB1MwaXm7T5SJCtjyONrmZXwRHUulLfxsmQAROWakpUJ3N7EzbJpA2LnroABbHPOvUVde
OmHzdTKHKJbe5VTQE+g8s3xP1nk7XoWZRWzQbPzqaQwlkX4mV5925qq+hLljH8FAQpbgiAMNFuVO
cNP1uC717//+MtQpm0xEgmIR0o1DUxK8Htg+0uI4cKPXlB0R+ETwdMWVXEXlo5uAShssPCfpsLXg
B1DMRm95v4G4MAR/ABp4gbT/jiIhwQwVu7LKeirWjkOoFH4koNQSwN33ydIX68vHMqR3TNz/8uV2
ZTdkOZTsiKRS4YLNugWFV7r4qYtTW2+m7zPQYECPqPzYLaIjG8cNbHtHI0Bj37JiyWtHi7EpLnnV
UWjprsSXIduOcHYrqtMf86a0Cb5lkwCT8pNzeeV9xXX8vD7cHuHK+cQiq6lLxkiqxSlnABbmFRdX
jVzgTqn0XjtLssDKA2qIBVfCkWvzSs655kFcIjQfMxINpQPa843608UJgUk1i8IYM6Wd1wryg5Qc
vHmDz4BPGE3opYjDTQhsMD03606bcVIqlmJPNltGN6cxKfgdjupRG5CQ6oOF/t2r5Q30eC0AZrOs
cWXaBqDEkmWkxD51QG8OUfY5460AfQExPIt0AO1dLUSl2hl9C1zJ6CAEgOjF13UNL6qKahwxuw8k
hYNPgVqdWrzbuzLESg0l/4EcFVJw4eU0jdIO1Cm8qjuAwQsBnaK9hqlo9LnfI4t420KlFQnSM6Ci
i8NEvfCWobeeYCp14ZN5k23Jc4r9JlvdioTf18H5RtEWwipYNIzRurmbvMgbLZDEQ1A/zbMnW3A9
i9epIR/7mHxxr4nflCvv6cWsrwwuwr4BtefIxGwfuQLtyZ3gFBitYpixBkK5U+IHwsw8FWxGP16g
whTmCLdOT+Del6XKoTnQQ6vNTK/Q/c+9ovLt9m0X61PQY2Vndf7hrmus/PDpMBAUuS7h1bYHetS9
WW+j6EXGYw9OvmCHy4nZHFnTRcO6UdpCrBUK1dKXa+Vdmd1oMPv2LJBxsCNveoodyo4aHslkj8mo
uSKxtdtnV3rh+KzOIlSFTfQkVh8sMrzGwhlLju9dYB9pt9xnnTUui9NXwy4vH3kNqotoEEnkk/RB
UGoB0MJfMjqOZBHklXzdav/R4SYq8htXtBQ9tUUKVhS1uR7EuV5CttKV4hByAkiIUNa5ZcJpmaK3
0yDI0Trc+d8PeKdLMSuQafVuHEASyU4TuumoZRN4fnZ4kYOL+eQ0vMd98adnOUZHawwgVz8I3oUU
ABGezi1rTv/5iU++DPgCQo8RD9i+b3yAkOZs4G+MOhaSUxTFBjk7utwQtw5abpnq5lCVOkt7hxW8
Pr/mtW2/w4fRQPCKti9YiqykhfhTVTdy0DSIGtCcMCoX4MYrW1+kvtaQqWV40BzvCE8IiplZRGeU
xJDBzvH68AwUzfWT6btmLdhpZdA73+/Dw5IISS1wArZlexG1ZYt2k26afOHFYRyhmTSYo9uR6dGf
z7lPVhR4z5YURMdno73E/mfYurqPhXWXZjI66nxJZJ6xEKaFwL68O29cF25XNvkrLqYTMHNrPZho
S4bBQidi+kndU8B0Jqd2FUVsAF8z/kufIsIEyhYnMmQFgK9n5nLRKtOgL2EyrP9qeCxSYTwQRs9j
bMFPCzmrUlfWMYquEYj7VCKFWJSeD4ijRdMvaw/nO0/3NdHUK8GMmdvNwFy3M+UcNTxwB1vPEie1
hAoLGLya2ge64BCaHn5k4ZUvtrnwCZCtlLYnlc/j8CFlmrjfmH5rGzFoprJDxhEavusiYOtNxM/P
INnlQ0tSubOPqCvKlFtbEe4+nGw9fY9TzBdGjFGYdgTxfmie41kqUL3CHZLjWtBFViCD6wYbTFeW
erkWYAk+qO3vLI7UyYeHBeosTH61E3kSYTApplQGXuZH+H965C58RIhii5Eu3NooEM8WGprdCAc8
J8y3NMNwvdm6j6KvVUkAPaSMTvWwGd39SDDEN2tHK6hkzt3A+5xdmpIHBJ5G2vH9S8iw4cTbAnWI
45Qc2kWYfmDyJr3vinDOFIdi/4O4LygeI9YTrDWps3wfrluaD2UH5cD6S/4u1MPTH3h43/Ai7ycx
N8dAag4EKWCbG6t6yVayhJOm0NUAadbsRcF/uflFVxMdk/f88IES28gwNh3/6YhvRgFHxYhOEz8T
KVejQDSfnf7Ss3F4cyS6AeY6XEMtNND42dXDdoDZiEnraYh33HKx9XSmHiQ/1NRoI7fB4ytLKe8w
ke8CVV/TaWMeEKAPRUGvix3E99sKXVI1xXBu9LIcdTZmTn9joKnXBvmrGnhsaCtaZT4hpapKxtdp
l8mc9Jebz8kzpkR9ix5OAOzXR2HzDeEcj2C64H23y7Cb5sl957smn2PosVp/2vfDNr+CEv1QeAwK
quT0gkhMWcaTt1BjOobtH2ykvvcclLqoiVFEPdOjVALs8jet7v/QDRivJ5wLfs3UksRrUgn+fSJT
2fgYROWU/QtU3WlWs8+Ppd19aRoLAQ+juP1Ax8Mr7GyMkwDd6aZPWqi0VrkvRMTBzfWOAErIbfIm
0fi/kTfcqN/1Xp+WLLA5TLqoflpHOdws+ECrLEUAthopLeWvXNexNUFUmaN2w2bfh9YCB4AyRTzt
jf0UMO8JfgxgHQ1UNKK07icXxt2CZM3xyHkm6X4k44nGQuZN9lJtV/YDsOfvpn9dLTtK4NVCYz5i
M1yV+Ze3xsqHShfbj9BLaHUE+dHRqXQcs8yLayRHGWqfHhZmKinHs0cqmX+cgVEK8TgtYI0qjuvI
HCn/xfQ/syHEwtb7mCoiTX7xdcP+4U62Y390eHzL5Hl4x/zcixDY4JKrXdQmObN+eaS7KBvLOj7b
UasT1LJB+Xnpcs1qLjN6+VNOV1kTDnDKS4YwtossLsQQ/5+dtR7yubxn4ez5k7AOFWrwi4l8/PxB
I4baIjuiWGWF6VVY0b9wWatU60foeA8sgYPVDcOXIK9hvPtgTnwuIbvEnkkHIMf/gX9UXiyoVzC8
NxA/DmqUUnoP4B4cSYGK0hKbw64/aFXeD7ekz4xPEZ8pBoYCowHkSU0gx67TiJQfWaCFTkUUt9Ch
TRoFhNiaGyqc4m8qjkuR9V7ppSsMcKuyefe3XJTBD7JU25cFAVxBIBBBh3Rkv3FrtgXQHfXw0hZn
/MLluAvjcLwUdQdjETm+MbH7tg47VZX6e/25aahD4l+ivBZBF8wopTziqKOZz2G+AjBefIypFYT5
uQ6xM4X2v3DLsdwGY1UvpXgL6cmMyAMAlCTeUNEv0Ab7JIW6dCYxfhZk56sN+fOJgAMEs6eR/R/e
MwpcwJgPfwraB5QA6X/W6JhdpIa6SVpCkUYPBQFc+v+AS9fEzC6M7XaXqpGP4uAzMmUTOW70Kjox
CbaqREM4JAXUOl99GHmLdQzNcWbLq9K/Vs1n3F40ysmlRoYtfxcDRotNephrPWQXifI8ztrN1Ef2
kZihiWWH4SMh0C47DMV/fkyPvi0A1WDFeOif/BwNGCKvxN6j6GmAPpmUiTsNIBxB+PkVDDcNtJ5j
DSXJv8Ti6YwulZD1PHKZS7yjnhg+Imo2lOQcbc/sRY7jtWkFNScBfXjEB7dURuU3A4dy/wDkCvof
ZibZo8SLkc2FXStqViV3YkHCFRbfkIZ0HzjP32pugCUsVJ4oNCdyIa3jIyj4toG1oamYqgMRUiuW
LmemjyJaiHTVH2PGDsQfKZqLaloh7Srn4GZ9qD4OxtyQ9k3NBQ58y4IeEe0pINS8dJVZOjyTWlbe
wMl+0nbaMpKv+DWQwLRLRgGT82s1gwR291KQyLU0GGZIYKGnUrwwFA0MKtrZgeFYR2uvJ2x9TTIv
6rUCgcrXnOwywtkcHohBL+alAl8hB/cl8jCQVLbkPWicia/FVcKVjCCawgs0VaSXBSyiNGraI9OJ
v77vGMrLHuF6le6D5Pqd8KJvDQPt34J2c20h2e7cEP7kFOpLoo9BD+S4w1qYipfcvi0GwU7EcGwK
etUF9tZA3UH3qWfwgbwj0AXJMwOA7LZax7AA3K8qaz/VGvwOcBloWrwfMPuCQHstpQioV2qIpoFc
306OM+kJyJHnTgw/HR/ECls54amwZw8bZsGr9zUEqHWP8m/heNXH9q3E+8IPjDNHK2a/U+VpZEwg
Y4fEk4aiVG7QmxlmqGj/cJBj4pDyUrYsgLtz3fc9mGqxA154F/8n/uYZngcJ8CyK6wnUXTDCB9xB
tEqf6gcrVKUq2+Jd/FR4jx5j4kawb8CoDXypjBmPsozzBANqFATroL0FrWROzpQRQe+qcGCVtKdk
d05r+1LXTtTpS70diPA+w75OjeGxqef0RmRWFmYhJMCtx0og8rLW9H4YQAIT6gcNf2IG4BWk1BoP
iMawmnvUKe8y/Bqet1zFIjRywz7rA54N7l+9HQ3VZsVFP/j2P/UrMDK68OMdjCLdT7V2X4RUAlEz
ZCS+SNt8kI3GqaEvf1BWK/Eo7wEXCA2/fTKEdHWWYklpYX/VA56yKYjl2SfSPAzyfMWsMNp780KY
DXlwwFDpcWBL29hCkoa4hqMxT19apjOt+soiuWVRnB3hBDH8Lkx0ToMxqVj6Ept8PhGEDjuD0Fq4
Er9hDIvIZqgjr37Iv49uudanAhN8bVMH93Rf82Lwk3CviAwsWbMygSDstoR0/4VumjIv32EOtZ1i
VmGoMq1PMqsCXnIgqcpSIJoGSolsflOmEQXX8+ESGepf8Vc9IxjdaEozCm1AyLfY6Lzjnm2NhsTR
qQcX6MmO/N4uuLPHGd8QutS1oj5hs9DBOkS3RjAFSnaKP4qOIZ4ajmugLX3yR+0VjcmXeIv4Sfn9
v7DUdA2ujrNEuCkYSpRQnAUHxEGsycsT0Av4ejJnILBpiZnJV/61HFmEo9521BjcYk/pnRRua5qf
8x9E79xe6NgDZM1xFEiNFUzA6sp+eET+Lr6tb5qcOA31vJdj4auWaf9K2rx2O30TSfxOZ2zqkkHB
fbNE7O6Ev33V2FZAe+ZGlHPtNnqiCxJU11+P0UgQLTXWFRkYTQlMrLYY0tuLfo7DHu1jNPnAARRz
dIOUUjlIvb8QD1gN9kCZAFJ6xb9dRJbDFJGCxOBVzknK74YXmtgSzWd4a5OqNA9dTuRxqS0qM/3i
MjoZIaIjXfjGgJ556o1PTioYAFMie/d1g9Bv0jYmIE5xODZ9fwlDv1gXJGv7DiGG6ZZaCNtdtGrb
UmQK41zBUtnYJMbTxBLSKH+bdQ055np0N03Di8OKmExjgIblI7yaPri/v+VClKDH0BdWgmqySzDF
lERVkH2csmlbPI2bT1Jo9xNMXnGPj1ZdPxZkuaGmmh0/c9t+8Uvowawc/TWs0RA1QTxD1HRbItiK
fC6SoUzqiM1Udd69qH6wGu6KUdwgeNLpfetWBgp7drz+s7xuyOvR/NJEuAiRGGD0y9wXJtHy3Ze0
fOmTPKANUUEPgvMiDPQj2s5WcEjAyvQawdKDkBc9/0ZlgTk+IQrTF/2rIklkQ41U5Y55hDNa83oO
pqTy76gVnCFapmDy9+CF6l/qNoDSz/vaPauTtjE9RG/L5W043C8793fsqi9zEDTySbWH0J3wIqFs
Wv8gwSCGoTkELz9hz2T9maHDHfs7S7DOmKk1yGiQOhJFbbBOh6S6eZp/spV+3DdqjczORUcTEtzg
s55iI9ftNuyWVBoH+GgGQ23xLNSosId1qA8CO4eIsXztDIImS8DUIo2c+5A5Iar8CvOk/6DyMzdA
WiopNqY2fYp/i2ZS5e2xutP9mjZnC5AO7aSvCj5gh0aluzBQtV/IqerPeaDDW49LCPyhsrnNr21N
lJDTXTWGRZs44oM9YrvZZpspvLa9tQVlN/xtjoZAyncKtQC67RQh+kZ0V0OoRN9sJk//ldWEsl4z
Ub1p/KVhCPCFLlOIbATOOaigctHV6U4n+4yKMMKFckXQmmD5WBYy6OutEAc600FmPURa3JTtZcgX
YiD0v/wRQ0eoigbkrxMJXkR3CrwAdiedKlSZl8MQ3ujbr269V1lKeoCPTKMksQrZV3spqbTGO1Yf
WBqonfEJgFtBxvHAb7jlN1pTHXuIqGQYU5oXfK7x7KxK9v1wZSPqNOq6UAko+t5EFWs4KqT3gz9N
Ul7JOcahw8zhu5VIgdWjTmLt79sAUaeUGsXEvECbhXLlN7mrJ1gJ5Jo+NBdHDvnOKqkBGIq5SHsv
vpCjUvWr4ozIoD7oIkgLFEzqaxg2CYLhbbogmTLauB7BVZ0KqqdJEv8BlrsGO4EZijnQ+xXMgDzD
KN6NOZZXMCH4EfoVMp4eSrbptKYVUdZhxSw2cCbwDEbzlgaEYf3nM6jy85KPhCSQcETjTeyjpX9q
DQ6Tjy0XlIJPPlRDe1VWdro/RsdL7Q2SUxN7IjlErrml9emPQzeFj4l0oHhF9j9mS68/tqQBAPG0
/h8He9FGkOh0oiuw1Tsnet+Y+ldWIZab5gRi6Pk0z32u89FFZU0AxFXNLHht2pQ0Jgb+zRCf+FII
E2Yk5IHe2SMCkYzdFhab/lbI9Plie1iC2Y44M5DGLR6uWsgY4ZJTI8pF5F8LCPRcVzYc3/OKsrJx
ayKzwvUjcXjhSS5LZFo3O7etK61oAF61X6Q7LFXzEKnbYPuzAkRed7lB2jRK8HIW1jl2IJlKPYJ0
/JVaonXffqY5BhBP8L3baRpRxs4r7H16FWdotKNJc7TxBxcWRbrLbPz2yUgi1W7Qw6faimKZaJBs
HNWWaJ7erkNuyc2dFSZRtQHATbvfYWrrcc7HkHG9RiI+g7tekfNkFtoGIV5JSGrp1TeasoVQv5OZ
8xVhXEHc3NUsHoz27MXf+QgdD6pJ1YB8Ly0YSwQwHGmpIVkFybN5t+vlZEqgrPX3ctecpeVifayp
nrSky1prjAkXdQiRTIhnkPqCL5+1Ba4z6TYgZdonQsa0sAMMjbZoKyG28PmWJksjXUHEA8esUVUZ
IlsB4uSkzkqjiMthg+FNzW1QhXeVBGURiF5yVeNx7QNldP4kS5MtD2UzGqji6JORhLyCNBlsyPrZ
NbEEhSF0nohQu6LTxFz6mNSWvStk4GQNGpdTfGDEVv2sKLH1mH2m+XXcFtnrdgXeMfowwp6kHXyU
rMEc89C+f3sWAAoNlGd4ZoNTlNS/bU0xH21BZQaqSQQsvrerKdpxfZoHsSO2pQ6gVbhBQC2nkKwA
bI90xEkSKIiRoUPP91GOP/eQ/ZQ9SFvPP+NoyDHrcovkBIJ8qV9KtPb5NLqgz9cL3OlE9pffMgD9
cXXnOqh6e0yZDZuFyVYzRmvPWGmQjMHdTPiaf55qxzucXcvqpn7za9mLiR+ycIPdEhfb56HqQNxr
6LJWEwyyBBk48x6Kbe/LW6ARBdlaJl0CMPBRQ+o9hYq+XytksdUQYJe0W2/I9VyEnllnFKaYCwGr
70AjNsxD69xhQu2D0qAzvEKtofjUz1CamFW9t/k0XvdotKXMrZ4zZ14qU391MlcAUsxibMGVKbJC
jGKKfWJGlYolKZgHIPnpytU3DiXV8bDcOPvhzIiRVeq9hwUUapbSLPiraih/JOpr+kUM0v0yUkTm
AaSKnCJZhEl9Zn0EBfQXIigsyCZKJiZZcmQWhlmY6A+Pa1lqMzHPgUBb2hgSHCGo3ldzlSYGaa0t
5odT/RQwATP+VC8IY2UIcY7bOOQ3j8+7Cn8rmjUU+TWU3hm1Z+orofkAHUMP6A60UrUjScIsJi3N
I+bphBZJw/6y2sGjeT0H9gvKIaAOggJF0Kv9lWJWz+qzXfsouR8OlY5fc089+3R6lznZytZMNPfI
rTU1jK0LfNlTFXrnmTbTL9i541zze8RLgf2PszMetV0hRSgJZiiiQXVbzPUD7rSzmxA6laFe1VJc
ur3VKZWpj37qPs6v7gL0ziKJPbq2IR02lYZQak/fntJqk7wrgjpmaKoXcAHwZLAON00aDgxbCG7t
VzTOkAXEVG3ydcZInRyrQWFg+cgyPD8rTS6Sb8BGZLRBBRB3TQuMGln4UHDTB3uIBdDTIcvg1E3C
XeYt7H3o16ZFDtI2dls/IaEM6H48QXhrbVUjnSitB1N3VSgeQlXMbZvlS5+zqsDlEGzAs4KlSfnp
qUDGO3I4OgYdrf1Otd/e0H5/GcQ4lW/Pmin7jOO0KO6huG1xyuJLnOqefHeg2eN9D6dqNLgR1t71
t8zTHdoC2V3VgYm6Mm0Q9GUnTHxPm3NqjyJ4tpYNkQrJSc5gIIKWaZRe+tQfxPFf5+BLg7vifqbL
yA1mRuqtk/eVZEwcUfbecIuDSFkH8vfvtDoYf6NMYYiL1FYmCSp+PJML2vLEEhwz6jqN6/3bUkkz
NAwtv2I6I5/SRDqMHKcFIXTEMHGWN+PShu7cbRsHdVBYP3PYfhxbPFGIkmmCC7Hlf+X2YXm3bZd/
/S1SnZo2rdolXhQxAXVQ4o45k/dlf/Edk66y3ihrvz3Y1yDk+PHokB71mzfNSzH5fdHaC/gaUmNL
LYq9eP8uBy0zNHOb+XG0zhxtFopGviUicgm6zAB6pJ0itpvQoqbt98Q2rtWU71Bqjvi9lkKcJIEa
mI8GU2OWC4qTIW1DR0iMtEv3TKhXghOXhIbm1kRlbLJje5hHy35qrWGGhsB0iG8yWYZr632dGXE9
h5LVEWM8uZ23KSetpNr5eoFngDagRPMVHPEXuQSMXjYV8KFUdN2cdRTRv50EuYYboJWWgTGiF8Vk
jEgdIM6tUgpiQJab924midlfSz1G+Ox5SOBMsTz8GMEgkEBxv4/AdslI/eVQ2As6BiRd5wtWlopZ
qk9AoqbFUkRzF01PV4DkOdTNeg/YKXwvhkHpm/1O4RWZy8Ee/w0iJTc29Atu+K0BIkb0z2u+t/xi
t6ZDPcY7P8wlvXG0onptZLKte/yYdSD/H+Uq8N59r00WqYTxtRXFbE2+z+Na+vDajg3coqFZ7M76
VNoHAkx3NvBTRQB27kLGmpLJsBUX7IsPvU3NMOry9Mo2ByTm9f1Fk2Wdch3K+ex4FRKUnOcnX7XT
5nFnu+peEzCJnj7Ava2WMqzzJ/EUbcUvgFVBH0Afipk8hrP/Va3U4Q6RprcD5ust79mXT/slF69i
LcxZd+CKJ+oBGmOuCtHv8tIwWahrD8HmG8hkmY4Y36BiegO8RVFv7auuz7R5VnBcUjAx6vEBb9Hj
rCNTpQBOaIS6TPX9oe44CWn3ctSwgTFuzuUlq1ztmgxVzdkCe3Ix+R4fWIHhyipG5TKkuCjsnlys
MedpDylgbBcOVecZjkJt+b4tjQLqilZFxxUbFJ0ip3lznbW+lP8MMmtzhejs0Ejm1PUkhWBN1cCp
iUHUh741lFsKJ5SSwQ51uitwCkyL2oYryBuOhT3sgASp1zJZmrVOe5SHu8a7VQJXRlQGQnxq8H8w
vXOdjV1d6pOI8P+W3+RdK+I41lEr0wMGzpT/uKtEKeVFHawRP9Z1xKb6MO1bgHH7Agx9k8xXI93q
XhjNr9ziuKto2rgGph8ABWMZlO+iiKD8rFU6594ec8ONtxeB+NeQ0NgYrbFrv/vPUkZLN/rU+yiO
AFDmvjyPu6275Pro7TV+M882MjJntAsqUXG0NqmJSLrRyCyUNs2NqczNelXWU0/oEexfepUkwG2X
gKfL4KEQ99Z++wepPIIVvmFFwOCbA7pIFg87/9PjveVyEPMjEXOn3bwN0gjBd6tpH6AJm/9RMbZL
gGvnBHt9Y6LcSWsYkONOthjKZ+OYx/PomqnbpMbGqDBQXQVoaNJ1hpdq3+YYoUwiefLWlJOMOlm9
Xt3gOMNuNmX0Bwv186fOKl7Q4AlxucsW3MAZoSgcVwAGWv88Oobf4R8X4LIxjNQXC56hkhz/v8vU
oBhU7oGV3f594TpsByx9nbRYoA0SnvomHJqtb4R0uYDG9OU2FW/ZzCZ33wd9B/8bMBMRVMe6bBiB
zCfSWq+307y2JCRmVInK+ukyOcshmx/atFK2c8DKaDZA+twpk9FoMO0OGz6Iymz2/G8kSpLA2318
Q7Wc72eXykNMZ2ePds18YjHiNyWu1D0cazOHaLvlZrrXhkdiAwBhfeSYxm74Kyi5eK68si5DTrWq
fgRJrepmAmkG/BgjFIt6MfUaHK+sm2qkHQGlDhLjAeCFSM36q2OkkYllRgde7jkgbDdTdWCjr9NR
ONAqg5ZCfbQxMsiTbEyfQqcv+nIdTcnO0R0DBMXJvyonHrsqRWh9LTo2xaUrb4M5goT1SEJhIwPX
JGcGRq6NnVW6KDlTtCpNBSmjJYa1YWV4iKMFHK8Bb4XFxMpMLyVWa8qak+hk7+FWH43AMYMTXYde
VzmOm0abKq/3a6qcWVFvJHhnjQjCnzFY4GFHjNGXrjwsfgUfM4JdHdxm7YWQAfC+JM8tblV13UTE
DPsMEC16uaAU3T3qfaRttNHLbEwDMXB4eq3ewg8XfCoFVThpazirl4tRvcMnxnLpin6d3m0DbrZF
8HFFDRdDeShQdV5nyC/pS6dLUhhDGCInD0YDSQb10zo/bglVj322XlM8IeBNvItpq1zBJWOad1oW
zT7CVR7xOve9aoZApJarcXLi0cECpPCoRJluWAkmyBBXMrsOxm1IKEh8p2PtW0NaW1RopM6KXCXY
HGcssfwc4jVQlhw7nwRsgiPZagXaDTdSQ44iadgEgSlu++PtA9+4YZl1J5/epYTwiYCOlcaja+2d
TrcpARO98ltgImEHVgFPhtuzPsdY1Ns1OpL7CsQRxq8cAe4yX/pJBeYsHX1ny+1B94TrDoPEUDaK
7zLjjXc10pNxnYujxwyJlyheQ83RY0Zkh6DTla5Lk1MN5lb6qHXVJ4C+X+o8urDvjsyasX4pHRbh
exl8RlRHYveEhO9b1eDsk+xlx+TQDsIfImK+ADBq7+mwpevHQVOhp70PvELdZpjg1fCYXo61wI/C
VSIjjuBDq+i1D/F1OMOiqgqFzQPaIMU8TzDN07ol6zPRrohqBn3kyt1owF7XqCq0CLp3DQ7226xC
LjgosMqco29Jld1MnGdRhSrAonWKyuXs734jadKmjlUIZ05wUrBI+dcSyeqk1rTD+veYXSAs52ph
hKjiICv3gftfcCcbRvzjvWwRnRrq/bWOdRtcqhnW6ZaAsK7T3BH3imX6DG2kzwPjJCIjriNJ7DlE
gLnPFl/V9CDHJcHI1SqnNk12lZIivMS+xAPCVQzT/ghZwOIYrRTvaviXQlGQfuOI8suUn6+mq50R
d8OFXBcHNXKkiqdkqGPOcVYPD7dYw4/venl8RFaq9he15o1vxF78qhRbNQkVqi5O5CmF6PrvfwVJ
mRI3taxRvwFrbuKE9aIafTuAca9JNyGCKLLNiWCW0lSg+uurca4BBNtUTRhLSzTw5YhiGBtnyFv9
DoEzQIXAktn2eC1XdLiHjSXJup6aCZZAmDmyGCogFZADGg3VeeA9BIxSr6SkGjnlI1lOS5G8aA/Y
IZMeWm8Zbs0ZCpssheSzxMCWucQc9XptVbvy1tkuyJ9fTMMuvMPH18JB0of/JESI6f38QU3BSQUq
gtFhOy5dK+UasFzI/xEhm8+tdWZbhXMgOxQNLCLxRd3o1HkcVVdlGwEhYp37PMDTw+zvqfbaSz1c
twa09LEj0f4VL7zSnt770ig/RoCrjOPS1sZeDYpS/5dCIhLMmi1aqSilTHQ/zS0zFIBEaxF4S70Z
MHeeNRJRxn4gkWW0O3EO4d0nXNdD41LwnfV/pDwYfVejlJUNwwBGPvze5ZKutfSVA4va5RsVX56g
x3R/EpvpomHZx/nJUYgJKrmYFavPGClv8ArPV3JZvOwVberbgNVSHrtpk7Med4SSkE4RqROT5LJz
4jQ9uQaYYJgYqddPPjw0VslbmVApF5/DOHMH4vWBjK3PMNfU6sXz156NmbaYQ8cy/Iezmr3LDaYk
rvEwo5aidekyXWOrngvsfUG5Nld6SjFkfuJoaPDygStCYCsyssosvb8pjSX/nfnDfdpUrgHCpW0e
7prLKGQLMuVeaVF83qYNtQc1TplUjhF2/rPNzH3PC8iBH9I34jU2nsJtKhBIW5N0oC4sATh8ubAc
T5dXB38/K0VMNaRAwdLB91CalnGIz2PAVq7YnQZan0cqDhEJNJvuy1LLjXHV7zk4vEYfNJiM+Igz
l+ISwc4rqEY7b/YjV2ZDvVq4FT6img6P8hRtA2KNzXKEgtaiZC25ve0jR1YUYEReNm1oJAzaJkNg
N/m5P4XEIM5An2Ia9WcsjPSRRVfFcFd4an5OPp7VVfdGg7JKt9DobO7P8fvmFWaPo9UGPPErIG3w
Sa7xY/qP9LbNtQe4DC3JEJ5OhxAxIhNDs6wgPEd70nMSXBFaRxyLytFzgCmfLEPgafO7W7uILWcz
bfpsQyLVAPsw1wOevd+pHIN1XnR1qbLuoMCuJ2lBrQXxSOU40ehqQwRUOqqJU0kb2xKblQSvPUN3
aeR+hspI5aErac3qRg9Efp+tBYS3DygMmfLIENHeWBGM/PKj8AqwZxg+q1OZomRYFp5C5tHJc4SH
N3bFQMxnw32AdK3lFiHwsmU3p7uJhZaIKwA7AMTMKgys/I8g3fxC00h/J7B9P1CkmDxZx0NXrWkV
LAAvNYka8jnlZRtnVj37lEfI/E/y1y0SFanJNB7oJLQN8M7ergWxVkW3kbRTU94z7qMujQev0/Vo
EtVG0LQ1AoxORsLGVTLLakyJj5r6DB3Dzn2fvJ6F8GaFGav/0JbzHProM1xUOk5KxE2msnKCKZbG
FGb06FQOrF/TN5HeSj6qv8liYeUqYSnogNZgumjuDc/W7OsZO26SC02WEjR7sB4KEGxDH9Pc80Ra
xQ97C9tcuBOHf6E7aSj06RcfxLaQM1YGKx9ndEWcCyPib7Ig7+iALKpIE5646EHvqIG5JJ9GP3wQ
1TmP5QVY46uMXIHEnwVjIz+R8Dr/0PtQ/nfluVreC2AAPfG12RNxUWYy/+/1+5qsvRE1SsBGi/NI
GkTTDEKTVbqFLrRvM7D4uPkJL6tRPegUowLfFZsa33jdc8fZ4Eos1iR+IxktJAxcHYz7UP7S861S
W+dZfcKNq0URxBVkBhJHhkMUeLtMLU6LCVLNnjDPqbF+LmmLz/cSuSkulGVX24GUybXq7g4jkqs8
ZEBXJBhWuhmrfw/s2IQYGUNwFTlAxTP+U/PmxmNKXidaEfxgAYCLjiFrHoJH1NiLdeu9Zy2RZR5U
KS1Oe9kG/mjjR3hi1UNqYVA5+TE2KY1akB6EC2Kf+xytvJVe+sIgSEmjHIbSHHD77nYQqk6hrpEC
3p2jmvr7W9DCGpYWqoiGbipCDfWoppZ8kroO33HGE+CfAzgFqaP5UC30Z7Z/BgLdo0AsxUU2fPIO
IsK04fJCJm4S4fxH9emNmjrOD2dRoAxJZHOATkXKq9dLVhfaLosiKfRJ7VvHI3g8t9faGRDEa3j7
8qR7ceD9p44Jd5paHtuw7/Tq8QevT+bcuxR0tVsEN+/GXbcw89Hf/8PWBuHkrMqK+ztKZDnVggTI
ety0+OGWHLTGTHpdl3mpYLqtsXTiGrOvkGceE5hcHrt6GLu1NjYQ1XtShkX9tiJb6H9tjj808k0A
ozpavzEpeJlXEVesGdiCQaqcVxlYLtXH50TUqe4+S9aX9dw3R8rpQeew8lImKbZ14YS4Lvep1Ko4
BOIwOSk3Psr+we2z1jN0qDwWbzvMCOgZmj1M8PTOzmg6pOVWJhQGgLNZhoyJFHwrWgH8GPztVZHr
wI9Bmo8/omGhA4teh7zVgYcyw1h2921h8JKOw0sCuscZGYMeYOKU3thdFr+CekIy5n5nR5jrUbpP
Eahft9SGIjrZ1z3WdNfjCm53drk1p+ni4KB0xEDoriLTvYJK3CiXt+oBdpr37l/xu2Dq8tiSPpMk
RSfTivXXuvVje3dmRTHEmptBnutGrRT4pcAC4EtRj+J4Pu2uKzAGJKYxUgl+K9rAdR25s03aZ9+8
38Ri0TA1blmRFyo9vK3qrHAQeP6zikaDsSxoKo0YjNlKhpMW4zT+/H4O73IKSuNEmFhteJAPsbqS
1xUaWXOoOFMCQeEwIMOxS1r2LWUMverRwXIKhS3XSZrqGRRixtTuhAHXLh190+CaAMPg2vMEkSEw
9To7Y/GYFeHzWKIKU/FiTUasHYVDyi0EdqoXtXvNo1TR2cyZjXZ2TajEPQ6EcmRlS92OuYk5qUJn
ixkjbkfhOBGTvCkgm2Yjp6eW/LVn4YPklEa4p7cDvNFAr7b95w4OgVnob3aV3ukHMxbIb0jv90SD
KIBUTBGji50bUJ7m0/aIkbJliNTOry2k8gPplT0PKV9OlRr1b0eIXkL06AWXejrsScTb68b+tpVb
fcVvlvjCFnujRlMCRpYCqPFyUQFI6vIjEXEakwf3KUsJWjlJtorMP1177yvmAjk4WEp5njIg1B6D
JK58/iblSdzFb53B/lPNucTHT9rpXu03Q5FaPHMmji9mQzPtSpLY+WT2k+/bkPafNavtP2eUwcy7
dnMOKYQkViEDioXxVv9yWaRmqMjkq54KqDXBG2EiR5wRPnXe0YG9/Mg+/S5DIT5QZWKCPffYOmzP
ycyBsQXvKxU4bLc6ITw3Z4JXuNSBTF+U3HkU43TtsluWRc+mxnjA4o4ZScwuCVwp7u2Hn1R6LmH4
aVO0qHx8SkJX4um8JhmNT9CQDX21lcKlmQh5D7rDYFb/NjMRNTOCgRWUFU5Czp8H+y/OdSTGI2kq
ojR38/i8dwVVzd8PJ5M/x51Xj69Ad1wpQo8MBrDWNSIHO0KRYfWQ5qJUicJFHLxJ+QjHeshoYVx4
ites9BSiHSS21szpRoQa08W3NpYtug81rAwPViSaQfTehLRRZ8Qm+V890AoWmq61e5tWE1Z2pUeS
H0l+Jl2QsfPwaq3+IE6/ZN8F/EObnWKL0DR+vPwwR6v0hQunLccEmEUWCSKQPfzaI5yz6P+byDfq
ut5Zv0PwTzVWCgXyyGqjzjd/B/LbPGWZtjCFb8MWNmUzn3GAXS7CHeKoEFreCVzi1+fTq+Z7Bbx7
a4vuAvObqPZCyRsGRXDb+rGNZ36icKryKs14JUutaKGSVio/mgLy9qjXsG4pYxBRJrY/8CUzb40r
E1sexVMmh6gddd/cVIe1PRpJUUL7hMGkKE37xBwaoEQO5bY7kOpHBMNe8RUGu/hSphxhRqVZuSrC
F0eCPvih4EwA09lN6QqcdLwldimVvcli7Z4jDsW50UVPSQytbUNxnBvavwuTWur3+tTWPZdk03u1
5v3cs6ayWwJEavGetg9gnjCcwAMaEVrCeTrLZV14xmjo+Fx6WJV8Rw1dEsOpY8ff/h18UZ2z7dnx
Gdha7V1rOm7iKg1ZhqgXVUCkdrOS85Dwq0m9tYmpPQL+sF6wAmF8GJ4JEkdr/TVxvRZMH2kCg26U
kqgcOXaj/83od1FPyzQX17etyJfszbRChoplF65bp4BVmg1jLkpRR4At/9RyoWe2AD1GxbZ1yWRD
9UIFzlnAXBjRV5t7keUyQOCQ8vmxSnhXMDBIK246CCAQKDpJrSnAPiGYGNv3beO0izg3Vms5uoUV
LAlCmhF5keNNwY87B4Az5ZA+2ya71ppFVKS5sCT++TDtgNRZLpIKQ4riewRXaUYk7hKcRXwYgoA0
rYCztsdbzd8jIP0Kf/oZ8tsR8ZUqJDeyzcard7eEYzrb0bpvIZY4kRYsbDnX8g+pm8EPeHL7jjGx
BDraBMJKcyTh7v1VKRVYMFsT2sWCZhJjj8Ye10Rm7xFeV4J/IL1oZIWZrKCFfylK4xoz7uJvWWRv
EGCGpnaYfheJ8f7YIzik05xpJI/Lm6HW13FCNiQEyONzrZS9dmPHyYcLGPLF2lhhpYvLOyyARHzS
jLNY0zL/kKF+dnY/46cdth2Gfjz8+CAsgx1j3LmP7eOHqiB90tYPKPm7h7kSZ4BW29fWrDWk5d8v
HS4eenNrYw9WlpuhtNOn4TyO9jRIU5qam3rGt96Uubjhva6p3QahYF8teWxbrugNzDrUdYh3p8Rn
bPwwUIN6m7pp5PZFILWDQV74ceBSw1OpwY0cpQf0OPPlccPs7JHe2+AlDKGlJxcG+LgdCiXGqXiw
agUuUfLCwiVfWPLiUlbVYmdVvhKBazsnJDvPsbzst7DGPt/PS4sE3draR7S1QGkrYK8imYcJ8Aul
dttM2VtbrEsxQyM2gMYWKS0EX41oaG58I6xyR3htxKv1yR5o8+dN1I6ljKi5Nmr0NGrbLwlam1VR
H5A0wLWI1W9H/L4/gOWUpkzdYvTCEtW0a+hrf9ahaymwXWZkMTuCDXXUfxdWqe1cJmnyojSx+hWA
QY+6cPwPBLksllMBLLnhYzCoO8P8cX0+TbGrPSckmFkXhZDsZvCxFfkESLbrdkPxqieAFzsaeQ4b
vWN8HFcY5Q0vyA8B+9AcIuvBwZ4xcZ8mhCHn4n5GXGsHLZiN0ctZ7dj7ibibiI5uDC+PF07Evi5u
3hqCaVjyUsPgLh2hW3oDLMT5lQxHNLVLQQDCSsLsdkjF+OEXcNdKgjdqYPQBwQdssn7CXfqxoDrW
8HvbKYYf7ZD/m9Y0EblnzSZZt+wkbFB+zOGF8xgvLboNoTunfStn9MTVd/8pO70xU2SHDSuuPzHb
qm+2LTjemJyrT9887aTlLVLm2PTxLmMD37Kd/IYMhM2wDhpDCwDX57Iixa7rPcNAOi07wHhEOWKF
DvC1CmapsVrpgW9JxIOcu83S45Bj3BWXgLzxtr9DJrELL9uK3EFuemoYeG3yn4w44t63VrxBtPNe
31sVSQPQ824OTcMYRWaqcspGDhUMGyhlbj1q+tETKtq+0+vJq7UqaHYdS+DWzywBUlxt24WTkSu7
2sfpfmUI/ml3IeFs7zE2/YGYRJ4PDH2vgOTlivuQw1Ur9vdpBSXAJVcKj1WmTxtuyuQSxEdyOVI1
hirmRB89UYwy1VxTnml9ChmBLgQ0Ex0vcr4FDGU/9DhEhsl6/MOyu7fD4t7Xtx1bu+R2KLHo1ECX
7pCVxK5UgZpkmndAKLS5BLEG4Ju1qrSsg7EWslvdrDV3umCsb8KEF/1WHHijyhxpnBAb05avxl9g
R8LeLtVK+LmgucTze/OS+K0ra292IGYFYFtShnUknUCQGigw7//HXKAmxy+eczWz0prW/KzQ5INb
UNNy+4k3vURc/DGr8h7isOy0nD/XBTZ2aM0nkaf+pJcHqLA4vshYSS9RbDRhO2N+YMjNneKALT+5
QFVVmK1kUkJ+Nr6hPk6EOX61I08UM2GCZsjI5WIbVsdK0x7z1F4s/3ZEMGzg2Nm/fRLd68Od0P3V
1oh2pGZxsv/w/VTfepML0ssD6aJqQ1pYer7IAwRBFaRHIAXSZ2T1D/Gl6XcW3tTlne1nB3/TKHM9
6nA/em39/fzO2clxmV+Lo2QaUNopU+20Yci+pq5yR1Ea0avzLI4MJEX7aQ1CJVKDZbue1tVFJgF2
2c0EWNfzkoufQA46N/98tdgQ6bVX5oqs96BE6bWSDJkXMjleLTdgjaFC5l+dIY08acXxrFr1JcWA
IA75iZhVMO2g18Rm1RRN0BtbV2QWbeaacndjrgwo933Y+WIEDR8QHKrCFtRaoDSuhdU0h/fwh95s
Dnaz7SPyWkNQ8MF+eswvsbaqxuAWkVgWWgNVw5uQ5PEC2II6/uNsT+lsjnEIKR2+Ck4UO8XkExPy
2pt/n2SMaejb/ysxDLsKQJnKGpZ5BPgJADq+B567/k5ZXGSY9teRzaA0pfrVWkg+qaioDXtKKdXd
sQZOoowudda9W/MNWnCxDuWB79e6ZnJjDpRincgOY75XWPMAB0blzR0EIdCvedrDkdQgnIMkmhan
evcVCx7uF/7HFSdZJvQaUK0C3GUTKEIR5SX65Ubqt+Fke2/bpsp5MyX5XpjqGxrm4Xn8H9Moifoz
2nysaRs7RylXzEm3A3xzolBgv60GVu5UocuqCreUlw3Z4Z8+ogElIHKd2BwciYaOhzzit8FWPqSg
pKGMqRX10ilbVfsgvb+7slCSZuOccomSMDtZfwJ6wKsTkhYzfjb0jHcgrCmGk/sYupl3O2+Sf4Fd
S2ScSMmBsBB9Gj/tljv30XGNP5xStesdldt0eLv9quQY97JRshEUaCSBL/SlvAVhJ5Btzlxs1/lj
kxjMKIRyQvkA/nc1gAJWw/KSJyOmACE7imZcTKkEpPMcSXixHsryWVkj5WNx0fetDNBYwKnErIro
9051SbqTkHbPcyZOJ2MWcl7Jt34R4Ejh0R/q3hyYexsn9/gd84rGH+WjXKAiTf8PzAKTkvGZ9fSz
n0dwmFEJ3DcwJpc0z04ZEhtv0q/l7usmJrfp1F05QRoi4K0Nj4WvJu/ypeuat+Jrd1kV5SJCISTE
Kj4pZnqYBOTu/lli7G8zCgzysaLIqc7Du4sds4dY0vY5KC3OB6o67AkUCGI1vjgASXVkMq8zFQPD
v6/+nnmuKc16/VTrx6Fva2D959T0BgaPLncTqemOSRxRrZsSlEnYqAnHJB2OaP2eTwQxXdDJnCrM
VG8iph5BX8dMZDjV9PKstr3S7uS8WeKAzLr4JeBC01nRqziI/7XC/yuT1ozMxO4lGWwc5/OVlMfK
2sJ7T6rGWCVN2CVwQ8jB7d5bNeMW8n12ySirqLaNMj42NMvyWRqMW2DkFwEapAW4hXYJu6JOChOq
9Ro2GtvtOYrvKGc/kTOEtEPqhJYgzYsdNGXF1xKQ/+Y3k04RF6HQXijtuDIw97rkoNXVBMh4dq9Y
C3G8IZmAfpRR8ZEmQC/K8cLexQ59sfB1bDFsmcaWvZbiPiaU+6vHTEERdL11oHXfM35F1LBDfJQ8
3+NLyUJoVSJmyEcbqNhBf1qpkeYbUeNbfXzOllLT/ARpuyJ7UQaSr2tSp/NxpRUVBzdGYjmVsxyo
/OqVt3VjmEpI6fvRXKZ4BVFNWENLCDwzgVXA1+l5sV951dcvzpfDqk390EO3DOkCbSgibXfrF4T3
93CJYfmTXYhwWmHL+QAQww2c+NDTMr8YB0/YMPeSH2iCBxs86yS+ZW7ULH7R/s7L5SCg6kOtAdhm
hyO4Jypcihwtckg4YFKnCxg2WHeT36v+4zZ6pNw9epJJo+XvSePWEKN82szrGDosRDKeVu+x+6Gi
Z4KByUtLUKSY47xrWPmm3TPW+jamvmg7sKKQGGCG0ATGBWF8dVk4AytV/ZLwjk6Kamzkxztwrhur
lE8l4SdWlriOQX+oDSnThm23tJMXVdZbT0hKonn/84Ld2mDhfRM4er3hZhxKXQDiN3J2SYQhyAi+
qqoMSbjpG+E+ew5POdEv5+raI5YFkzsgLve0u3AqXMFcqm8LEvrAAjTba4NshGyQzES/kSM0H83i
V78kFew+UGc5bkucvSwXY2VooUebWbjPNlzciM8Jb1XolFvJUJKYvEimR6CnesD/XRTiu8rzV+uJ
lbAGTKamDdPpVnzAEfSBB39lDwZ9JiJFxDmfshakqcs0zZq1pCetldbJL6cCyJNAJHAi0LgQedZW
JWoWV+v0lqbHGy56Fp6Xua8Kviff067e8gkZ7l+fFVAxLaMUtvehZ8boBPHExnW8l32oh3wR5/S4
7hx8QP57NHIOJH0zOitw4KzbUA8LPbErIOSzEmn+1g6F6dZfl3uxNFZRHVRBXWhLdf4XvRGQgS7/
dZQopxfRRGLqasp2HTRwR9X31jffBsyzBOsEgzpXJYZhq1hrxtsHxjc3qhCJ3P5TBMsAryEd+bNX
i4E/rPrSBGkppECA2n62OWQ0Ln17rkC9jCJvaQFjscNkoJdcPJfz948WOG4bwBmVfoLmToEIxC/o
5Nl/sHCZuycQVUmVN1AeSu1t8l71kvyk38cPfXhqgmCzL3vvBkik+dwyy2v1UUYnfvxzcJ4NtoF9
wqsIzBtzI2TEWq1/UBMisU5Qj4HhSy8htkY+8w9ZzQPIrc3I/W2ZaPIGL3eRnVHF5h5uIio6VZFZ
CplyLbBp4tkrFdF0FVAECFcQr+QrUqYBcXUNx5IRqZ+eA2m6t5krrfxAGYyGFa9d/7WLqZiXcPo8
fc6DMaH3v5uEB4EkLufGtFA8JodB3vhleh1MHrnfRxuxIiT8WslvuUHcIsBi25Bt+ol5ZgjDQj6w
iijCJl9mwpZoN7M/+k5F+4adl71MwnhlzU96C5IvsG5KVR708C8uTGcQ5uiVIkEy84wCfYuVcX0D
YI8flnkfzeliAL84RxOcuIRV2WneXx8XRJBRIHA4RTQgdYD4j0W2wXhKXFyVIXzjO2Z4Vr25Cb7a
7ZntpWzOf/iKG0TFuTNWtOr2a5Q81PYTgw99aj+NZfLDszebtMcmG5rnFCgxpkFImi/qBL5ogD8P
Ica13jJhxStU6LxaczQIj1z0+MrEKJlQ1heqPHwlRXsv4giVdksSwGY7EvwcSkuImlOu+/sPmlgk
KXqG3Lum+E8Kr7c9bxUnJD84WoRX+Y49yQxsDZRUpHeCD9jbezis3V3YJ5lOaeAvqLQz4XS3HqXD
GC79gJIlOBcp32DuKSJK6wZYab6oMQ2n2Fm84udpgcjY09ba7oftDATneSoe+uWYxVLFqlHTqjz0
G5lD5Tt/qAzMaQME58l3ZGFeIGfem1k/1QcYAhwtC4FnRkK1gXLYXg2mSnyLZ+MyLOD00Px1/Zxg
ElAhmc+q1FrZlGoFFvMmH/mpMf0K7+MVaj9GnuPA8WBwqrcSo6l2FYJwQi7d0Yi5n16F5dIl6vKn
9+a0S8TQclc2orvOa8oyK8wQJums8Df7Dqn7VvyVqxKATd/yrkmvoy0KlKHtLExPrE+FnIrH3h0V
uUtDr7w1UvWVkD/iaBwTGDO3EGy14BvhuuYM4GlGZcL/nADq3BvUsnXOX3+OWn3UmrGBYMmTDekO
QDVgxWSkPZ/aiOcRvQKvRs+Cz+ufM5SBgXf0aSd6rB0PfRZls1b/AzBRplMkaWBJyMVoehhpbBGa
dday1Im2sz6aquR372ngWsYksQ04XInpbG5h+r/GQzX/ixSGv/l4hxkOgmJ0VxrMtiG0o4cpFZWU
AbpAV9Q2Lq6wBVkUkKi9IeZ7BMxXn3qWgYo9e8bYoppl1jFU8tL2/VapnBBH/zdpcCRAx5KsidKs
t6KLWcYLkQeABOH0oUUtnVVgUzkioC7PeHvdAfAOGYXAJXeXNBINkLUfAP1m82BUP+oI/baQM/44
TjNDiPH/YkK/71wxOdxk2xPxGmQCZhGCYx6dyjpISGPq6Xz9cWbW6YQYSdSVHajCCKSi26VU+/H7
PIEmzmOEWTFwddJ9wwZCaDVpgzSjtmW6xGTYJkWM6WXSrPrPQbCa0JPimYBPOapmWTYPHIv85l56
AWth26oQJJMuMCexuhhp2ObIBdXFS1rzkbSlbmEW2tcIQKYRahoHGDKDnDwnIu5xkP7vfQHOJB37
0nTEn9zDeDpNwu8ukbir5JcfDHeiUGcyqADTOPoU3HSV4ATmFmuYvYqBt6vnbc8C3VTGC9rQhIul
yfYcTT78oJkp1AaZYP8nHW5EICgm+CrzBN0yopYILC9J1/SrTR+t4ymyKDkOhwv+Rits9G4g4gWy
YUOWYfkX9hOziuexd7ZYSXdCH9mtbwhouBqysvSoH837/H7OEXtuL2BBBsJONXJub+4/YsHsGPwX
l4lQIc/HJ+vxuzS3uoNLgl/SVtdCJwB8sSwKeHlQV+yKDa35jQSYY6tPxKYnUW8Xl6EFgNBYqvkO
2YEZN3EP8XKMuZxS+UAYir2cp7ZQFYRNE7xrLhh3N0c7+rYUS/CUbJQCgusiSMuRLRefLsoXQ96G
wzD0kCJxPbeSKdLvrGvkw/HBHZIXfMJ8dJakXTdp/ACh0Br/VE3KbSwyHB4nP1xUBb8gxZlSvS/+
gUXXaDY8aTF5mCnnNWBY56docxmPabJ6SA21oBlmvG0ORULrqLAZOCTz6sLxEvp3iyxK8eU3ELqc
3fhY91FpmdTU1eyLebulhCUUce2jGhUj4hgJ2OiG2GunKD0JpkBTJ/0vmYCaE+xg9UxN/2M1O8Pd
ujrYQeGJHCo4wxiwbDuOcNJo3a+m0SMA4ohHVKo6TAaCvw84MxSvH8j65+rTphnjR5nH0glbyS+y
ghTpWly+b7yI/9PVH9lazEuwvVuDL6oyXf6zHA3RbHeUrrkGwqI9ViouJTh2XxVg+sQo0U69sRFU
XekdOoUfGZLn1w5yJwrtA2zCCLfia6Qt5RH3Z6/adZKqd2ExEjrVKc7cH5nj6I2CH2yxcrGHrCwH
B/ExKkk9Bhcmiv2lwS3bMBGXoCV/BXugH1lPnDA9tzhis9SHS1blxT6p+x54R4FXWWP4kvwjCphw
0mMmeGPQyp/l45YyIT6ZfBgb/3q5BEhoNksynpMD8OQfZn1lrcVWeiwN/d53Fqq32atWTAUGxyHE
avAJEzt09lt12YwuwvBAH4Du+zrHyDR7q0RKiTq70Oe2DslHcU6iI9UJYWNlYnz3FeS8lDQ9a2oN
VUhOPsNh0ljtD/51wVdwPoo887/1jGG8EvR2e474grxKIvmKpKFktIM/J7UMay+CxJKfw4gNSaZA
hlY3RDVWK52flXsIsUhLs3Z4k3DdeR8TE/5RJiKHyT+jxjhqGFhXsxJ/nJDeku05JXGCIAYtHq87
Og6n9pgeSg8sSvEzTcl9cLniFHyeu58Tv1+G0h4WJYiYuva/lQ4fMm8iY/u0igaLPmYxMZ6MyhxR
4P0BYqfZntTD8T1mmqCnZmCPa36+J5FsGfAyDWa1++m1RMBESjw35tfqV/x2OLJY/lYyQF2k7DAC
MCSmD8UINVr1qyvokbUjenWfnjy+KiFUoZM3gWzr7HB1zXOrd5LxVhnJO7Yyf7/z36ED8ck0G4+A
hljVj89VQZmkGCyOc45Dg6bguS9QhR3sShFo2UPPGRsrJDpZDoIJMF6GlmpW7Bsy22xGRGBI4zUg
J23HLivsB+a0udGO74scqRJtfMhYXyllai5Ohw6oWYoefK7099iPR7kMyK8EF7YmxFbRPsVu/ImD
jWyzOM8C2v9JzfUV+OpREr097kcF0NKYF5lrRNd/7UZ/WVxGmg7icgHYnKioYl7vubGeYiNS+25a
CXKCDxFll9/DtVsI+JEB2ezExfir5hhi+doeQzpeQ4f1bZiehsV3lFqZow0NniVW/Gv7p0OUzM26
Fa/zORBkTKmgZG3G8Q5qy2BWPLOdvaKOaTHCaRtmyYlBMBjY2wir+KcW9jzhh6/yQd5H7Si5GHjh
qWoTMwrOoRbEnaU5Z7m5IB87aIaiU5zRwxZgXrUYjv8fntRi0RTG6EdCkIiPQE9jhmZIGmB/eB3X
YnDJjX2rKsA1LI3aG+Z+WnEjP7beTbAPgvoUN9+wM9vn4zfO5dyahPQIs1upu9+TnTfy+BXad1X1
VuAPWrhyRKo+z0ehdk9ctjqZVMp8AqV0mMbBz1Us/tSq/6xbtj6BrgkKtIPc8xV4cWa6Q5Rva6bM
e+ih69qVtvibmJUiZeU6iAuRtXl4E32anLUk3d8bculCwq5AvtKjQ4NAi8x8+pg2zUrlkkgSfEIX
N0Eb13y5HIxHtuRAxgP/bwfuJtatv1lWVDk15sessVV2lMZWMVQxmvPtDU0ZbN8y6cBIdzxSANcr
LJgyHoUUA2rjvkQ/nNDhknU2Ujik9r+NJvfztgla+7CxCwHhwXvUTS8kEZCOCVINuUhz45II4/7z
VhsFIXgAfaJ6oIhsN7mUXb08e5+doy6S9L5JEkepp/3rFYHCj1H3sjRSTgmzSafwCJxqI3sVTZhV
dSo3e+GwOWKZJrHXNfY2wJM1KhHg9DN33KqAFKAyhisG1qxJ8ni5Jt9Wer0eLBg/fDWT3+qxOEYA
PLbL1tGIrKe5l1NBpwXSL33sHQ9+hS5WX5KAc7Bb1yOkj2unYlPQJS3jKMIGHqlD/oPkTNsFGqi9
jVWWUyrETIcLrt8T+mWt0P9ijBAFj22O+VklNCEHljNzKoq6BuyXVVPPRlBI/fovfMMFs0SjS/11
6E3WehhuTvM9/Zo2jMDjwPt0K0w/93VWze9NrrZYqGP0reYri7Pmvfu9gga27ukMPSuDG23X8JfE
+Iq+JXIXAUUFAdHL0Zv/M2uG0Ecekw39o9rP0VRuxeVyZ1bfdMG9qDb7WvGsVdq65HydAnH4FxS/
EgVJ36rANkBedUSI+ck3WPYEt5Nc1E7tfKtMNA0UeLOlyu5xTt+d1UJtmdSytZkBtzq2PCqvKXdy
yIFyqVSkA0DEalUmor2Bahdxml9YU2CZoToz29pQYo0v72xLIfpHQsBtHYpX91mnFlE33fxkBuQp
IpzUsNbDb+RZEm9YZiYvSycs/bNyQwMv6t2nhNebPXeHoGuWtLtm3OLUsFD0oTv6smuyM1v1rybn
7BhdJvQ85UxUVt0ui2uREe9p83kGkqx7kx1sv6Rx8tz1n2pI02AVKkeWbFmVSCM+/2K7w8IvUbdO
nqGT9FZJNEqgK8AQdRyWQW65c+9QlfvGmOhTbYtiB+vQyftdpflD/orwB4qeREPVrN0YhAbYUvNi
jbCzUFDqXYz1whQsHusWSMDh30JTrz4JaynH/gAVQ9oiFYOzmsnVqrPLBab8KKkBNh45OcFGHX6l
jqSv5AacivRTCDD38A+QxyRVYRxC1kgUtp+neWCNjjpBjuDap41WExgwH3N8aKiYZ+EiJ06ab/zN
dHyyJENI0coJQyi79bk2AxYSgwjatgkvEULQiTiMQn0/G50sVk5tQnIzxZZGsn4I2ph4b0TERXam
cj/6sIPik2x4b2jum9M4YuKR/8HiW79larMytjBmdUhQChtjza/SDU4Lfug6qEXHR2GC3WIojQWB
WWF4gxGkFRTd1BASxCy/7V/Qzh95UzKyvhotlnLrXLY/Q+hlR6i1JJvOFRVYXMYccxgIYGVz53pn
e8DHyLGnd7J5Mh6xjWpEn/2mgkeomuoqRLlOrFN9plZk6COQO5JgUlY20YLKmlcp10xx4+ftqIIG
QBHzHvhtBAaq/BuOOoNJ9jhMCZ+ypKoTPY1eT8Sl0qyDm+HgRM0R8m0D0XkL6wZ6mTiUlM+157JX
wCNl56t3qA7NVL9kFystd4dAmfFFTbY0hj/xXDZar9dunrALTSe7d6qow8XJh4RX2CSLko8Eyr4H
DZx8C2qCAqinbT6t7rlAK1Dk2KilGA89Nq1gww5LsIyr7yN32U/wbETx0Pz4s39gyM83MM9CkAji
Lj4RxMf02vM87/R1IzRcJKjFybfDi0sL15raFntYweEs5ggH5xPmhwlszpt+LuZds59uCAmakUyc
kJEysggaiWm3GkOkubJdy9J7IJ2HhqGgEm852SRUQfoUpPlF5sjzb2CTLBli7lN+VX+q8InWjL6T
UKjQ0pv/Jf1bHe7EV/IsS37SjVvjfW3WhyMLWqx89OjCDZhQoMNPsk0zQELNf6yFNqQxpeAwtf2e
60dgHaee18YrWX9pBz8RDE3WP8l/ED8rS+aDcqOYjN13WeJxmzs5v4whv2/zbY5u0RXBJUQTB8Mv
H/KtqpkpEQUgti68FserrOK1Kegv5Y2wbxFxua5wWyFeK6ztDJMlNmDsV5kOIvbBsvrs+o0aTpo8
CWPIRJOSLcK67kwKFlt3GczEIK/ZfGheSpvpLMjzUU9bV0SesBY8FMcgDdv7F2F45dq9ETnKxNi1
KvY71S2MA/GLshKL/bMjBtVVQ6bMv0T1M4+B+8mCWrIzu0012EyedId9ATt1P74zDuBmD4BeMUf8
EykqtggLYpy/i8VmdlU1eBmFXqWDtV701t2Z4pFmP/Zxze26uOKMzIItLv+1EqdkuK9CO0PVLIF9
FoMt+UwnR39OSBkkIUPdb0BYDq/wX25JmwIXsoEMlRyndOoTOYakzv1LDjLD1bGq057Zh4kCn+su
UTMl2AczzYLdsiG63cnp0pDroccJK6ohlm3bCYzIOQjhChwPUgB0xJ9tY1ZujkAJ7JDgA2fmJVlx
T+Pj69zDw+qtzjcRK1Z8L/oxFZ9AVpe1RG4qfSs+0VcJOliHuCPXaWkqAPMIElJGiYOPus0lSwrz
c937Scg8XwYyrqYhODo9EfGZbuY3aoHNtj63ig/nMNT1Twua6j4lf9ZSPro27eOeJGZcGOz6rtUo
OtdFOxREGsGcEjdti3ZoyDg3kU7lVHDwpy+ZGV4939BdbApIeSeJRY2nqJviVOjvrmM69+8+msG5
5Scpvz8HAgzM6vRsS7TmSa6EJUmTpz5Rv9eNHIlvaX74/cd3yV5SWYxEV/EbT9x67k2TtoiEdkLP
HqkTg42PSvCERZuhDqReSTwHlNcqtZUUM74vq3q2TVgOcoNLuCV1E1YlTZgHi9gzUlasTU1jRSBC
FtftHifRKoslE3FQf6XImDOYDPZMAprAexnMA/Ty0doRrTGDshWZvGVnTKj24SJQHFOvubJmqO46
Fwu0rvmCd3Eh6GcdW8epq4fqGJhxvne9aPiLDsxxWJwwd9XKiwlqxYxfGtf3izmxUlqucOmvaiIF
U//kA2p0plFqvNL3PzfZjfwur6MSPQBqzsSUH9Ok0REyVKUzitNp1mn5PHExm3UkD0LJKe71r+ip
9+9vyErNiXL71etgCjiDG3yEK5wg4M8trzJc0RuZJULUO2FdaiNpwZ53g7hvhUVWcLb+DeA/m1M8
ziDV0PtbJHvTY2R+HFNOUuof2uQ0ER/LairT/VWnrUkgQPUoax2XSfS4YA+cOVZ+0Ye6w11gS5mb
Ezkg5dKzizuqpXoKQKHBsRW9cKSYxqGo016eBN2R/1p/IpDLo72xvfpVlz/m65cu0o1HbUlQSKPm
NJRk6kLA0I1LoxUnM4gdkApSi0w5eJxbkYBJ6ihaMjcblIUDOZoAG6tfL6yzIksqVZx10L3Skplh
9OhGhBUU07NCtuY8atO6Tuto+z/EPPJnK+1jGFAU0oD8uxsa3hJVdgp1He9ExD0YwO82yMuW5NDO
DcEysnmcm0PORCo+MLY6+LmG5os9kY5yBmz+RGzbfE2GTmjh5nfzQdJI1e+nEkbAF1XGKlI6BQnc
P+Xgwbke9TEh7mdWhHmee9k6kOuVegLjWHa3VWPwNB04Y/fso9zfu9W4OJZ3X6Jmin78rfOky7gV
hv901K3d67TCT/wqOKHUYgnoWeuXpwxJIjyl4xP24GFNHwBx/+LQFNKJaV0+qJC9GOpejANdfhBl
rIxebbm8QKHl6RY1C4NMdZTH2sES4Yo8KffyH2idUkrvab3hoPgdCs5BBwF3Z2WIXqPKqpMQP0Nd
5U+cTTJZfSW1NS7KABwGyllvEwDw3Imdzmyg1gxrPUManNX6XGsYjCWbu1ghNkJDjDLJlG0yGqMT
lclLwFR2/umonKHINHDqsNUJtqqrRI3Ywj+IhhPUGYqTv5aMcbA+Oh1WdsUB1whAMUBzZJOOkEC6
MgwDk4O9CWq/KCb6EarcJyEWlg78dczz4IUr5NmMeh7IO3w5obLtmh5Qu6D5jutuazQlMzOtSajo
+yRLGMIQQxN7QgJdkvwjd1aqTnJGzBznEVm5Co+j8hmtxWFKEj3NH6NLiuTdY2lV06SKoLEaJElU
AC0UQ19hPN90RNXOGehcolBMoFRdUzl3SWs9KSiDynqfHjOu5IexGqd3nuypHqJN2fywbgY8/Nt2
yc5qb8x744VDPed9lgrrxlqDrGG0v57DaOl8AeFbCHxkYitu0a/CfFlAfmb0Z+eKAHVfceOWF+MM
QHnMokSkP/SRc9qPyMJNQ6yWev6LnZVDQMbQ7DdvdB3RBC/7uhmQGALqiU2T4Wf3ViydpuHRsldR
+QU58DkSy668QZI1Nxy6NUc3R5ofM2hjBoFHQAntGUpotXmx6aBUBfPmOqi1LdvLWW47QUZ9nuUL
86grPKS5tZXDdL+Egbd6jNagJTwwKCVPywP3lMl2UNYcAjrrhZxRFnpgGH9TneSYrErmzSE7oYFJ
5Q5gq3sL4N+DHXqeZ/PBqBA8kqiycRgA0YbpMy8oBG4+mjIjdHICcidvbathuolTN3nu1/7F3W9A
YuY6uFjCnAIGqP+L+JooLR6VGvgwcMWnig5a8T0sD7g48rABc6GlTDboiGN4wk8CzYxEFpm80BVR
a/xuGNf8MebpAuNxitvZjgXLLJC3NP6xtttlLgZFBNAVj+qvXbrYssTeNAOWr+KDtAGDksIx3CVw
Wt93ZND9x2jKKkv3rRBgqgZ2bnuHR7JeFwPcPzht/0VM9pehbsh7wJ7/AneI+y7TRYl3JifHcdc3
RwlbfGGCB2LSPQYcQ4HopBRV8w64OHI0nb1T8jiVGyIJTuU4Fk+2hx6obPtInPo1gIya2ZHPy2Un
9PGV7+2dG00RNYXasO5z6m0O8cwsDm1GDvMCeV/QXcDg9MKDyHvq3Y2ncR74jBOkm8zKOfPHA8j6
Txj1F0r0/rbGyM3nhOLthcOUc1PSfEHjReHVt/Dw+3KshyIrmr9HrDwWToZJD/Ib+iP+Ng1Xi9kV
QD7UJomyyBb/8GPgSAlFszqZ5UXkQEw6mxCd3jaXbFiv884aRu49tB98Vj1CnPZlAaxAItO91hhS
CtWcaPAM0uUNjpjFSHxXgokOlENW0lWsiHQAL9eQ0TP0xO7UdotSB3VDW6XDp4n0RBvlHm4sT39s
TbkUAv1AR2DZerc9JTDIDW0V1pWVrXO1/NqP7xg86qU8CU67MvpbMuo1/J3pFbBvmSmq0ywxgPix
EyUB5Fs6NLMaiXZa2Qn6VQrRvP42EuakGpE2DerTJv4c8Y1rAcY1RDI1n6RZcNn//gHsVyCNYCj0
k9lzMKxHVqndXKlFpK8IX0m/CU9dAJcDjMFj+h3Yiqfkbkz3EOKjMbNHkcjapTjuXEAR8ByItDU/
rSKyyqPDa90iMUtL9tjg/NYqgcUChIGd9tDrI5Y2FWWtMWGRGHaeMbJ+vfccyKB7d1NDmv/NLIx4
pI5mqZaQiwBs8jGN7Ns8L9Np0qg+uEzQZpEDflpaoGf2ujjhQ/d7i/Ev/W5MXiRb9iicsHcMvkiz
OD9qPHNjvkiWNf/9kWUyaqHRQYJnCQSOq29l8QU99xPDPI0MPL4OKCSviVSlZKrd+bUQN5tG4w7F
NmLQiPaCk6T/V3SB0Z0dgtH+/j+Q5w9RL6r249T78XcyVweeKtaCX5kvk2gJkaKeWuLfd4EOgBLi
m9FVeLMBxnv7XiNMIFTv4aFqC9mif4N4fiQFRser4VMSD+JszvhXN6QtabWtTLUbRGYaV1LOlcH2
yrFHRLN+ftOOpeacCynBQy4qJtTemb2sYjb53Besq8HyGivqQnPgBpnfAwLjj7wofzNU5wUJbllK
WcmOSAxtEXTWBtAifHPn2uAH+GbOjkvA2r7wKRttw4AMhOd66S4swcz1AzDeqpdItQu0Vb7URmo/
PN69Cpq0lT3Z9QQ5TvXMoDLuc9fVoAR0g8PT4iW6kYUFHQFMWZX9/+HFNV1tlgsAILzDqHrTMfFU
Qta5ZPXt+4PRU7skpt/vDGI8et7bLsKE/55ceJ+UC3mmuxO2Kz3D+DHDVJfHW4WurY3cnKGyRVE/
jAEOvXCeNP1XSj6Swf8OcLbrNMVgiIR9Ngolp+U1nHzV+dXNy8+/LGXWQPZSVyMlI1v9zmxZDRdo
D8N4FoYf1arvNyBCUgbvll1cr6oRVbiiYZbTrbffSa40x/qEjDxfAWeOW7Re7bJ3jTx1FCPWMHli
PuS0y6rC7s+30gY3aupimyxCpXJYYr/91jvbxv5JTVkdfR3S9KaSXcyjatsT5w/ECjvgThP2Zm79
7SSDAXqRayesEdtpT1KlAReaBizGErhGnYLekyzNvX57PtS6serrC2BWFWWRmHEH1OMEvXHxxuXH
ChJ6N1MwrKkw2oyhSz4TNHqFam3iSrKcoNZyfAWFyeocZidMEVjMwWoeNnO1evq1OHO85LLPCqXW
rYv82wyqxD1Iloo69/Bkux4N6BInjbfURwOtCnl9vwNyuULvcQFsDiE703iy65Qe125p8V35+JGc
8MJYaTVHnxNMgvABFfUm5tkOAiSetsfgxKDzuCk8WP9Db9M+S3HS326CsyvDWprlG3wNz3mIxTD1
IOIUivkuvvd0Rf2HtV5BL2a/pILoYK/cu3PALSpDsS6w83ecQlRIgaWDYvzfR1p1us/oVsSWJosX
04yKvyphCKuVM40HpB3W09Y/kEkcrSl78BqIWcGs+KvDu6gdQPHk8wZu2DwXDIVxtxf/pdGxjptC
7tL0pkA53JHuICnwWg8HnHGeY5xf1tICMOH7wbw6mdTi/SwWs9fMoujjHaG6oRPatx6AuuZuauvi
tMmbkOWZIVM0AkgJ9f0tJ1n9ob0C5aU6zqpLgderhrxSTnd93dKvg9Q+FJPgMJR6o2V3z+W0LFXo
hmdpADZ87fqVxdBVDCi27AHXee2uWURWtzASHGW8WSwRjFSkckoFTmiwQvWoGGtLp8LWeKkMrPXf
P2LC6IV4gVU/ETu5vgiRIyTMCpuPYy1m9E/3hS+GD8EgJYeMdpxv5j9VCPG8Cay8I3ubrz6/nHfW
R7kSRvee1nVIN4Ht7kjn6LVUlLgfXIjyiFaupxH0ermVv3tBlZOqwcG6e1jK8qx8qmVoIod3IMnx
+q9wIB/oKhBijGsDR9FH+rYwBYIeUyiRI/HJaaVMuh+6q9xHsOmAx3MMcQhYS1Ow0No+roGOLd9T
d4bax5hLl5x5pTR4IywDuaw+MxWdQvIb60o0Jre4yvJdXZ6l9AFb6mKt7eJUcnz+6EvJ6+bDQibx
VPmg6egPb9j4sgKQ2GeIVeL1vlP4VDBhauwQ9F+celxG/YhxyMXBB1TI/8tD6Y7JMf1OD6GHMM95
Zxuuvb3Whb21N17FLhmVU6o3RX8EIhUpXie5zYHgrYKH1lcpmQ8/mCsSNJoNf548It9vWmQN7298
k9Jhh1eG4w99gYeAURp8hyntsjzOEhoKno03DOHsmbzyFkxpXaa3GRMl6LS6SYOv3B3Qtoulb1Jq
XCo71vXy2q8dDTCkMlSzKtTb8zl/CVLvVIQ4BzhcWqxSQDdcVRDZyHnoymEaeZxadjJBpurDim3q
2L4XXGKaHTFAsa+Nw8flVFcUSgwZrNQswBAQt9wkIcgYNB7OhexxhgvYEVM4RASdP5ni+5bnGBdj
+u5IcSGlOuix6xu3X6tD8tawWpMRCoA03w13OqrP4yDeZUWF1KCkBOt01sWuEZiMZlKK2/J5TxoA
fn+rFOlBnWYnA97f1BOvYSILPM60AxNJGnUIvPscqySzbR00Zz2/ob/7zomX+jRdKD7bBm+EPRtO
/ZjdCuvufV84THs3cdhDBa3QYUNFC2OfyHmU3DmbzKZ15NwAQq/pfq8SmKxfgEt1p11B2jtwuyDk
73+FgSwpyDNzcj0tAF8+iCqMTbuEwiE86NKmqlkt3HrW3RiQpH+qEvhk2UayoLtEn5auGpv9Fymv
lHOcdaSK/ZrCtpxhFk11fZsVod+8R/zucLUSoJjIac49QPgP5aGK57YUoE50M6I1/jh26cLI07mk
w/6z/sRNVsC3syp8iUAsCPPoBCF2ALYBKNWk8OPYjheUHHLq8x7VcJXR3vzO9BokwE7prYDpCYMr
p7tIkEc+VrvurebVAJ4Raa40fcm9JuL84ggnlyaAFqS8mV1v6gFIAsO8f4rXE6dfzzsssJG7n8WG
tUM4CO1mmVfQtRgfN5HQz0InrUy56F8WXQ5WWvcdycLPKbwlSriw9wmInTTH4tCqDX7UU/RV0MV1
Qp1yxoHGiiCQeB0O4pAx1FV+yKwQt6ijTcKRpv6FCCtExVc1tBjwnTANGlLXFDsx7xUkG2MpPlkF
UcLz4zVKZzfKJgrCbLQQAJCIQKbN3vt1NM1W5N/rBk88qqKG1wmLFoVENNLsxx+Qc6Lbi5RlKjAw
f+BJvkQ10fMeNRwoIV6qOduzt2N6w5mp67GQDqLYUWj4PbQd6sKgnIt7RlWkthYZKUsBBGeykq4M
ecLa9iBFwpozlhJB+YQuESs6d+LFrDxwy6/OYmdL9tM1r4Uo+R3ezg7V9bpcp752HODVVKe4PVZe
EgTmF8AQtz8rqknFUWFSPT8pFEIoFOuBQVj6ysnbHvXUzXd6lKDqhPiWOGxFHXbBJ2ANhumBeLxQ
5A1v1Ii27F5qQghcIFl4ZxiJ3mwvm63PmUOU1ZSlW/eHWDyeixhig0nIO68Q3juKPqSFbzHhwCEz
oEcFRmepDGINYVhmKpkoCyYvGjfR0W541irGf6HNdMiB7P1MDTv5jaYuiXahd6KKR30my8Ee7Y7c
y6QcjO07lg0OzAsZnNidP0rCFScsOhy495q6at31LUqgf8Q83+TT8BQ78WZXGzmyb3kfEOWMnOQY
cnMFYb6Ckhte4WMgSvuODENIExwdCyMmSyBJ9+M5obTc3yvvoYtg+G7HBbBDH8oia4jKm9+agAGi
n7hV5FzGiJhXFZhdZIUnsvlSR1NWhO2bNMW6g8AaRTSwAznXme5aap+bs1qjnXtriXiAmUh6zVSS
EaP8KEfRrS7zke8GG+rGkm4GMDuroPwEVstFJ6/aOTyeP5sYg9oJTN7m6ESFdT62HuwEG5z4Xka1
aTXnlwLso2tPwhkCTzwlReqIUBY6ocF7Cil0PjmVlnYQVQEVUO7SacaTL6zrMI6Q8TD/vCRnESO/
x7sg3D0/4xYrWvH9weVD/L8vXDClWXTiNGQHRw2yoOXl2HVVdv9eiuyRBJQg4yEhr03gVOU5VfZh
liLsaZ3dyi/gUzH2awQ5NCA5pM+MwVm4iLnRXVRP/j8wIA9rUC/UvhdF1P0XMaFmVoE3MLgI19ml
qSWI01P9t0Pe0gj7hdUEDf9p4/+zCCaTs3Eem+7TZHC6vypYS+PWDN9RUtks5N5zozyVGnFkqUT+
otOvkl7+rRnrqk2crelysD82L3CKCQ3OeTX7aFPygnQc69wAgwBhI3g76DkApPFcb41I2fTUAEG0
/3/uMaBm/qiW7/XSghCW68/2w44pDcooyOZ6t/zzx36Ab1rRN+YRiByB7pwUahv5kpCGE1KYCKKm
DIh4TTO9eHmTlFX7xDrwJlq4Fb3sUqEdUtvKxAooiyNN6N5f5XZX+NNyzR78XBHjCj+g1bFz7Ept
t8astU6DIlbILuaJr5rXR1noo28dipxuWfE6uU3Fqos0idjQXrtPSVlABlhDbWgRTTQd+u5bprJd
yDzN0gfCcpxI+yE8fH3TGJBKe1xQ8Uy3OkRS3vCYg0MZIwkGrtVlEflasVnUBjp31Kz7agYzbH0Q
xnc2s7SmVgsjd6WFmJIgLYmbY6g5oJ5FJmlAT0rTnc1c8EGmTjfT39csDJTVdLSHE8Yy0FCPq2cE
G+UGDxhvjkfPm6cDnje2FVVvwSJOAcZbCuS+nHI1Lu2hB0RWsJxHppTonSJoxxaKT19W5lCtj+5g
OWAd40SizvQIwRgs67f9LJYhzDI/nbpJ5/lI4aTbgm0MlCEzMY4Y/bbgAekzhc0kvhAO1ZGBJL4y
15aZGBYdeRboGDWuMEqOH2u1asAIw6uMuKvETRVRmugH7SyjnSjOqb22qrpU1b6P2FD2T0Q5hWRS
VpjS96BuSzKlwZZv6ZjGSB8wtLWnjpuIRHZF2yzEMfL+tPsNf6e2Gv1mTNsmEMIDuUbUixTibjma
rLSzyCWA6dXqtUHfMV26XSImMgD93JthrG8f/eXETxfCieFh5AvZxYspWdsMtydb5Idffb7tHqTV
KDDyXIie/IWX9menEHSMn3HsfIDOofNDG6EZkqrBDVN+ykwP1v0Z2SWJ+JJn2JiIJOaamWE6HYBb
unA286VINgBjx9Cs1anOWWKApeaGOiE3GJuKzBGJh/NTGMng3M8ca9FTNVlUZh476ebEzfTUQHCh
9AxLJdFXniLCYBcSV0Y4CVt6gTnWIzBwD3IrX4FWLU2Ch5A5YV9d+kJdI20aCg+tqH97T4wWeJ4H
Wf6QSBapB9QRUGNUFbfLeHzk9GD2y5gM/U0yJSVb4HqL0t4myZqjHQh+9WoSYslApwIYkI+xAZuv
EREVHnFEXCJg7LLoeo5vtTxwA5J7QBECdhAh6hWwN0GC1kL3iMSWL5DJTXuUrWUGKhmO9cU7ijB1
JbNaWXbUlr/EXyQfX9ePoNgUZrDYpO+M4DFcO8Uhny9PUpaTZPpwTXMP7rKZrcg6FWSaNmwfZsrD
5woE0lXthf3RhBtqv3/hws5zM17GflNuLTnWeTuoQwBUW55pv2+Qq+ohPzNniigJyNpml/3nGD2H
7NpI+sB5/js85MlM2NIe6BQSmKhK0CWGntptpHVAcNMQrpA4OzXEDmPVDNejMICPKfs3ktJVmUH5
Bi62RL9N1T5G7jFVSKsRuGX/YOMRVkgnPIxajW8IypJc/S3HqJqIm3MIK1i7+jyKt9bzxN6MdWXc
rOEQ/I/beh7654uWC9NP+Tgfggx7bAViHV7xdprq/0cFuunph9/u7SA2hcVPKXurad/01dDAKhM4
Cz4Uo4q4x1W/gIG8D73CT56sGTi05GLZrfylFN5ifG/2baBgHNIPoiThiEZVKdzb/rk4oMC/wcmB
NkjBH5qPgSL/v5s9hwxp8x5zjYpyGFHMgzdBdbsNM1KpZNVuAmVtD2fg4lKExEYOIK6Y8XxHJtn7
JnDaGEdrOGOoe6CUTA0GHvO7VNa/lYtzaGQ7cjEBDeNX7oe4wKCNV29gWKxISyo+CjOuce/nua9E
4T8xOUMDOYDIJTG4bw31LsV1SpNhc2V7jpbcZT817sdAX+CuG81SHS2fG2n1CyTNt4nEmeT+evD8
GNfHSBypV9iOiOsYW7vCGfMfQH7TJ8RYFgKICZjOdmsddSZDTe1Aq5GAqDIA/7t6gzOm8oE1BrOc
JdP70GTwm5XtHtnwqFCMaqBpws57VOfwup2FBwgxjbNz2So4uzvBIKFy9hJaqMflpd20YZSCMLIo
V52VMSF0pCYeo6OFHp+HCWUzuflRSmPVghVmhxCRjJQVsqQgjd9pcMYiivsuxCIIN4ZmyyZS9lCz
r/9EPYJ27G7TMrdAMe+hj5VX3Ilwa0qazIpuMKnT8z3k1ispTJ1/a1RDO91vuUUwtVX/aeUtyQLp
b2DFnBrQ+dhsk1PpBmF6p1rmn3KAlF2NHGvSeA/Hd0uFHImcV1QPK5kcjayMFweYJPJFE3JOLNid
YDiD/R2pRxQa0y8Wd4g/+TGY96WA8u9m/r/u5R/6mBwJFyfcIC74oN9fc7IM6mGpQ8f/i/eSyJD1
b0Bc9MAIVhJSmvgnASm3gkDksfxdaxZzrYh1DtHvkd6SnBY6/+AUERzugAefe8CfizyW3asWBbjJ
riBqPzBJmmiDJyM7JP6Z/WjyLokQB+Uf9Y8I444hAKCS7giMTR+4g+1MlqznhYWV0uCOiB3BzQ0F
+QvkOvGjvv5vj/rYueRQ9NR4uAs6qyVAegU7jKWcN8ioCQPX1p1PTqXrGTwwQm46ZBrxJ78pG1+o
7h+PHE4HZCkdQIJw+2N+RLsvpPDrnPC3Fpkdy3r+Ujw8inCEo/JnNsuPfocyBYgR6X7qQdZe5D7p
eILNWe5lgV3cReyMKlsK+6AtYqaj0dz7mVZb3m+KRg1JU/1HQNZe5nGQwHfWDJvAzBas98vxlxx5
Sf8vH9evSkU9FpEiIY5St0c03b7IIsf5yTbWoyYX9dqejh99AYPjtUGK/yDBCAz2BseK/5ttJPj4
fIZtvuCBvtU9PbApvLkyI+kF2VLrP0b/iaVhaaioIw8TpEglK3pUnhUJxwnNPMa0wZeXawm1AR+y
6sjne0ACUXxwO5qUC95kYWqRLJkdECqtCfKfeOcVewfq2rUnYwgE6n+OKOMbVa23FGipSaULlmrF
V7LPChSmuWi/wXWCP8zVLM9NDWCnxa91qXOHVRcdt2VRIjzDgUdlzteeFwbk1hExGRbmRO2ltRHv
VWPDRmbJSHR6F752QzS+D2YG4LPCrvEwwKqxgylcFDHhnSUFQXUJ0fQswfOO1W1YbnlcJjF+yzlw
Hh5KAWbZO+08JAtLVzPEghAXIGaZdNYTz7PPovnkDC4zTTEcHXyyJo2IQ5N9jBdfPPcVeU6LqRnD
ODekX3iG0y2jr2NGWuPotNURww4p3Je83K92sYS1zA3icqT4FrdkW51eQa2XiN6e15zSnSmLbdIF
ynkl3DaISvGpj0WG+SpHBbLFv/uyj5/usWzlD8HaQC0k0sHcI7LabxJJ3GkLc+W2iHA7IIw1wX2p
cMa0M1nz0E+gRLQW65Wvp68wshltoVVJ+R4Do/W1gIy0iZybxg1Xlq/mISUzA1RFj2JOg9Ix2zgr
Ns3PXGcsAFuo4Iq2whXctubUhyyzIAv6s9UjbjynCFKSDm3N0LVnhX7rLhKzEOnxb1zzw/PnI7IT
5kbBOHw/PlNwczW4dLJ3n78PxPTxfEdT+QYhYdYc9vTpStMHE9p8+LMUB/hNW7kwGM2it4uJDCJy
RCLEGzah28J+XCWoQnVmESHFbocpLUiC81NHb/QJ9e+9YuuHguVBmbbMgzOeEGnvn8N0eGpBomoM
6DnptvF2LDLyhga2ftfI5496+jPZimZ8U+UchUOOvXtvVq2Tnh9DShIxf78FIxaxIBJm0F95EsQQ
SWiZCqQCaRDwlfaxAOkgam3yoHoGoarnfoGwB1apPofOWDmwFpzq7cjVHJFaDGUo5jEsi+6/0uri
grz7hw9xoAv/Y1gs1DTirX2DV6wh2f8M1h4yH84e0Hb1+bmu1Byhu7JHs7ZYv+m4JtdJSJDygilP
x6XLY86G4kELDI5uBtNWtHoTITKAjwlEfkPLm1HIrq0xqw0Zh90RodRNcy/JnN33ld2lwT0ct6M+
iAFZUamugtWdMBDqb2iH/z72iD6NhRQIZrZ8Haiu+fanqI2tARq9HHsTSjkYkvfws1vcL30tZFSU
CYx72hjEvDmXDxCGOU3AeYEB6AXJtY5sV7ovH79fgkPil7nDicvPeEM/hkNn6dncym8pVULytnMf
xfX76V1rjA64gZLp/pOZNZAmGQITDDQENQv3N5pAEVvRQRrLWU2+2UutJmvXNDzby79AtTkRob9m
cXIBVJ+BaVAqtwr5YYdJwlkQW/cdrhouTS1ljt2fanYzul/OhIOC14slLwiHnk4AvtM42wIove2P
6sLNJ/te2rGt5U24xjgjp/nNBWjbssvataBJA6lCK1F+viVlrSZDI31RBqHjhrBTM93aHu4ViaJw
oHCa3H9yVoeksh7G2JVEdczDuTWndlStEJeHFbnHZaX3Otubdym8iftau5NGZI0vAwq+Nu5+i8Hg
Q2xe7sx+H7orwauYstXAEqy4GqZ/sdteQc9ZmM5ZpSZo3Ri7kJdmBE+WT585/mzNV0VtjJFT70rG
7kkdZc/Gz2sKJVf1MjU12XUKpTobFDs3DEFkuigAajSYAXmLaTYGNgxFkx1lmsBRRt0wVXVEIr/o
F6UtC5jBJ1lQoTci1uPk9MWteMnXZVO7gEYWdqT4euasB3hiKYwzb8JXqeyiGJnguufBv+FwGkWn
d4uMu1xFosGdZB/wdkyD/5my2WkYfnAcTiP+IVlOqIN4jNWNNHT+aZcdLB2+QAed6IEwqmXWcSvB
NbwisgN6CWG476fw1tHjvaaIXq22ju/4oxvgsEJ+vJ2i1h0gd36gzyNZbt1T4vM6E/SKuxIOAWGq
7qJjblZUFdQBIkMd1XjY6/FDeyjhLcMQwqSM0ZnlByWYez/ZKqEGYCU0uDg8+wx5IZJNd1iakyQY
RdITNNrc63e3PyzVDkCbIROgHEnmhNC6cAxchl1E0gVyu4nVnJnOj6EI+N9GW+5VPUEvr6/yDBmP
KHdpfgclJMqwHZqhFKcQJ4nof5ZMdzfardyowempWOstzcF8i0/weq3AD9vkhur1F2OZlW6Fapjd
goiZ0nXM0rPFNTQUm9x4xx3QPSeg+qtbxXoTDHFRZHdlFk2Fx5e2ZZpXcc6Efyrlt4APg1hUSTEi
kTfnS05J7CBpg179ITKGIcb3cefQcormuGAbW0I/w9pTEGKHBI/B/u9+I3dBem6BRtaO6rd8fq50
KLGZvHyiEjTQGm4c4dyoU3NVQNAMzYnNrd1Xsh/Ws9vSB4vELHftdjQJH8GM8gspcif+KgKy8kaV
n6Z+1EdT27YEYFYGSETTx8kS+4h5CQeHyxHPDQvC+FV5lNuOvG1C4GT/21SyKp/+N7eHbUr2JQaI
CJGjH+2hRVR1URxH8DJVSNHzk8vrVwge6gMZ06dvsjZPlzjHDtLPJBPzsEmrodl1zDgT1CoO47yJ
zKoFzOpOSUnQ0WhQqF3GTnzQstCQv71F+PWlntn/LBwrwSCiYt0HbqEeQz8AMz+noa7EyHhEEG5+
nt4UnY3USytlY28GSeWERaiigyxNTtYl7DPY3iyl+WZmkNw2DEHOrUBPsiIp1UkGIPZEjA525h8p
F6BZAxoB+fefu1QQLVvf5oeLJzGTImMkch/zU3amDMtYqPBMjt0sux+9zLSiZHIePE/050cFxz8I
76UGJhXz7DQb4E51foABPAufHGW/D+9XtoP4mdVbNxbh0aYPjZK7HeGxNLNDwvyPk4EzTsgpp4sT
xaU/ajyxF0fA6eRXUtLxhM+ggrLu9BxnBu9ieAeA/tKTIWdPihqbkn2dC9PBc3fadfsPw73HKeQN
OmWVMN5wO+3HGB5kka6KMlblrzc+WtbjY8orO7OFGBE9MiMmDV31qWZZEVcJf8UB6AW0K0ZzVWFl
JRO3S/4fqPTgcmaO5Oo/AGHNPLpCPTyn9qBUPRnoyFVDxXdnvdmlWa0O0iKAdWPde6XccXNTysJN
8B8cCTYfTWPZWRhHlSBJbNZOnMlkMGIVWHaF+anRrUAd9tEe4NP88WNLCG/giWLothDw/sdoeX7A
y14RadIzIISWuq63FPPB3xeqFXk61gJRDdb4QbIi1meIrvmFB3eB72DOt5gIOR+wSNbw6hzeFxqI
MPaMxHHzOtXRdkqgsdTK6cXYcx44mYIk4GwbN6+CVbJELIEISm6xQn2x4QozSk8ZG+74L7qh86Xa
obfdLviPtNvzQS5iSb6ra4uSJEJafiEsVkT5XPjiWb4D6Vxw02sKeJEXW3rIqOc9r4hHrn1NjJGV
oHX9ZPobl5GkxPQDL828IPcKFGICE5yuOpTJX2joBlfxzixHe/lPMlRZwnNzg21JXNNmRoYG5/8O
EBm9ckulASGnfbT8frSTiT0rt2Ok3s9yqm39jBbALYsSuSjjiI6y127U9IcgBRQv1jZGz6qi1vx8
VcfqkjKWHBn/HtvdKYV0tx0gAhnug9pzs+v9G1Nr7NpknSQlv3CMi5pSqkhpX9V2c3j1WnVq1FiS
fs20RbwHc4Ln/un4lIW90USf6z5BmRHFc0FPFsBGofK6OOh4/fq06OltgyQtqzD7fohYoEzq1WSD
HcU+XmesMAISjXNJzS7Vsy/Nufq8C/lHEGnQvQWU+tuqWA17prdk5RWHMzGQ5HQ2oi7+x95cuiop
X37LHyuwqgulPn45VqAZoPS2bqlS/zQWmxDON7ql2cn3NYSMV4fe1p3BCR1s5X3dLKXkszjY9/eD
fwpRiuLRO20QpzLTssmY2Y9rgoZC3kyOafIdhDPapKR8V82mXhxBik9xkpfcySQUY2wVxDfbN8ZO
Fu+wsX6MV9SyBOxDAl39MeXyaQ++GMq3Um3TW5tUi7Ip0hnPrV1+Bzq7X/xk+7TQcHOnAxVcQdgf
zmfWElklDrMSct1UKJnoHmoJG1pi5DW0u+UH805lJeJDp4WK4Qamv/BLLpvj0e/PpvP1S45ph1uj
YmUFXI7RG3MkdF1IRPvVVOBOX8Q98JvzVXL/b5HNzWrc/TY+PXyAtwwfWJxauVw7gIc9SJhGPYdp
Gl/pg57SJQ+zG/ID+dioHQN5T3E/vuZ6wOxCgbfSbPeqY1oLD3PUyZg6H+abWvplt+FYLVr4Jm2T
etHKdhuhtQ48f6sK7h/5DgzUrGIjT5Dy94wgcxyw3YQrERErQi63DLhMGEIT1hQ1DFzFGL1JJw8X
lHutCC0LAsmiXDIfymd55or1Jk1imY6DZabfHcdJ4F96/iyqugX8z5xV5qdpLgQRuc0x3sQ1wG48
xY7BoOU7MyD7C2aD3IL9HI76UfIyzB4I65N/YGnBwZIgfgDI7iIzHGifOwQrOzwSjVa61P/iXP0g
Kv1xz4pG1/OE5Xsdyy7v9tVAP6BIP5i2KA4eDrcavkCY+y8cZAEOGZty7BeGvW/J39xVQADv7GOb
mjUtUKJ9wSWTVdGqLhmVhNA73kGbZRAMVJajluHs8T3IVOCNc06nORBVyV6eMyDO6B3CuKUu9jGB
L8lx59MsUXn+LZ0LsIl7fIlnz2drbfriZ06LDeUyMza0kg0PfTB4zNU6rSfENKLEXIQlXRm/NNUG
F7tWn+afebyWqmQmqd4nPSgMG8d5BgmXCeAJKz+X3KMZ7us9PMRM/SK4nXs1BdSUMLzJx1jHhLzb
+TiNsXj8lhfmJhTlKPsiQtkUraMVZs7Hx7auK1ecGncOvj/h5zyFQQDe1kR5sk+ZiqG9NUbLB8P4
xl9uBd8CHCDzQfvjYlWmCr6EprEybKOlRhWyYRpjFYv5ohgzW7BnZ5YyIgvFVSlQU2eZ+BKUrfHu
N9OE5e4fiWQa1p0LWZBwlSPsRIGUOaG/IPZLlGw45kbrLTNx/98eJxp10Dg5EZDEuZC6OtuL0fFR
nO4AXufHt+VjDRiJYBMnluiIPMJueokcdDZnIELw7cPllYNtmRp6vUehOHJlV5jKsQPcex/plOom
D7uqldZBJ0MkfPt9MnwCBx+XQ9Zk2wLzbFgDe49RNKRa3AKXi4MPYQ5SGqS3hHgLBpurITQYcW8Z
GiXCpc/dWO4MeFkJLTJf8gIe5BTQPMRRVfJB0Bm/banrh5Ag/hc1XscepIYMvtsEP5Ikd4lgqSv6
cUGsfjLzDI+g5oerha4WSar2nH0sttAKkz2ZDsh1KEBlN2U+LT9eTdO0YpIGFgQepJVLU13KApi1
uXdsvejcU2+JDqsag2CPGELjRbuZHZ+Lw6+cF+15fUOKb7kKz/+wGAVw8ULT4/6RAEZll5/gKrFZ
7270xkinDvghVoCWE+0NmWp3MWStZe1OuZWAc4PHjt2CE5H3lP1JASFymlqaIG+Y2FBpwwqPhQB6
99BEyuZ4k58d6ohOtwkpKllSzbQxB3xMQuCUeLe0pBCV28B/4Xl8Qv2Ifv0BfRhgsiiEejK9EU0G
9xW1Ow8KRwxhib/K/2FPB+w4eufSvRI8iROx0ILfVpLYElbDADriuAvgVzn4kOfMPKKejzDheU3A
weYK8y1sSxeSS940KQmkN6pcapF5E1P4z1Fms9Zp+GBH32DPTL7rV359ezZ83n0IEKaMQu+G/JA1
2ZHK2C0MCxz0wcBrRhm6swnmP7Fkz9R+gSjDiUaWTYu8Pd37jVNonq0BpBdGQQTAGmjuKkzplWt0
SRpnTGxN2KrOBroX3EbEhSQNlIoXcxVX+akHJhOqh6aRhnlCX6ZSEUzH16X7wnP7CgQKR11OeQ86
uE/+nCGpOeRmwKv0xzRasmL41ceCeEAKSbZ3Ufo83diOUz1yZBqF8or7+c/MoD8JV2YT/c7uW1gC
0/1uUw3QYo2rz1GXhTH+uYoJNSVp/+ys05Gk0Mn8auI75SUA+HNhsShJs0AIcnqriESSWZRBBOrz
hwhIBVKXM8l0rGZlyIDfBGBZYdrAyJbLQyZ4/7Wt48rv/w0RJfvzJVrNJ+AonK6xDgOP35CxE+qa
TKIIHt9VAyXPs58Ia24Rr9qrvoI7AXfxiZj/Zq21IK7dlUCLaqt5Z1lJ+iRYO8/aeQx7W8bCJ5it
MdsVXU5osys0y8PkckZX+GLyH3lyC+JUvQUFtdRttI1arxtd0sHk8aH5pZu7FcymKI+GbkQJnbXv
5dnZj4M9o6bLjRIoFm8Khi4Q5OQbN4V1u6/ri1uGxIcJRuW/ZamTNphE6ANZFY3hoeH+oN3zj/SO
bfFJV4DYP79pUBd1xgMS+ShVK44V4WTDS3N9uPKox07HFcjPsg2ogKW51KqbB/lkEZGPis3L35pR
SzHZfvRE26d0FhYjfh4AD/k7zAtGhddJMGrh8J8ShtvDq01sdko5TNOwv7vTC/Vsr6iPaeoGA39C
ue2OG1Tvt4C7mXWyq8CfaQKrDTbBX5cDYnFb+trKQtDJdqGPoaqDgizRqfOMAs7HGc2k1pZgj0Ng
+4Gj1gl1u/gMP4ojdRVsgKoW7zNxYrY5/gHsFMoc8OK2jGO6mp8tiMKK9lPYCzWa1/U/1x9fRpzg
242gFD0HbaHCvfo1o0RL0Q9BhMRcBmy3y+ECPTsmtpMo/JeuDbg1LOBa2cUxzHDdHHmSpgXbGm/6
LXD8g3lq/mpm1SyiirrntZ4Uv3r4K6pb2RXxde7jDrZEuUd/AVoaBFGXMuWDFJ+wD3RRYUvCt1sP
tOn8eMrd162fjDs4GP4vKnaf9friHsbX/8NCbCgQdAma1QEg/fF22bQnysECxqpLMFiSk9qMO8He
URQ1XQ9TrW+Ni/zlWrXeiKX1jbN1F2wAdkBRPUJ2QH5m50aCkONe80F/C6UyH4H6dDGu0NW2S6Mq
uA3Pj+PIfCcoAyctM1ZQf/REeNLWj9Xk1bjFWo9zqfVQ+aitwRmXpHd+H+4m6qIrljheDtPL5vbv
ccP9txQf3rJfR2X7oaJK2iY8xOcVPQ4jFzZb8UJQal4ypQ8AAU9iAAsmW6J/El58rft+wzEP3FkX
7rOyYm40T/SebkmdNvWvV6Mj1EzEnCneDHSZ1Cm00SF5Rov/MxMZk0b0GGyVkUWuEGS57thmxAC0
bPgVxbcdNsHT+0JAmmW4zNNpNkmitS75MN0kBZSMyPNVpdoUoY8IboE3HPI36y3FvyoxgVcf6/rf
QguxyHlF+ThX+xaz6tfu+ZzG6XgCTU+Y3V8argMLAIEDtOcu7WnDsg7djw/Gyt2fu/GUStRM4g90
jK1r+ZEtMQf7JgWFs1ZOq6apX9z5tMasZBm+9KOVfPezeoRSWI5cPqLNoqwG0TJyh9VGJHGEQLx5
jzbeSCuFobOOBnUqgX9bnqN8IJ7xz6GIaT/ot//Sv864A573VFlaXwv+WK8bcq5f1MuawOnFOCuP
epTl/dE+SfJPJp9+V+SJDQw/BYEWpmKnWXRlMtojT/6o43UyS6+rbwWqWgVAd8mOaMeGYnyZZood
ILNZBGI6fuuQ3Dczp7qaGNVW4e+Ro5KKDGXRNjvkAEc7nMGzxGKCX0XJZIOEfSwBZCLU9ms84rNN
owewCYwSq4CoJXbc8fEjYqrFt2MJadEAmIL0ncKNKra09e5rP3I+lb6ub+Cq/f7bJkqxY2EJjXP7
KA0+NDyIQUucJMGYC3lmWD9gIMt5CwuIJ69RtpsVH7oAOUWMPIQ7rEx2CfeJ+/K2AadO7o7SPtF3
5LQ2KyPNfMQ4ekRRDQD/rlaEMtBxkHUwDSUUVFR7yT/DW+vRDHY6JzANu03OXto4MTYxZrjm/fe1
iCbnNUeAjXxjoX3YsEhWiWrfNTjnZf+ys+oZ+hLezMMIWxWlvL2JWOm1g30xL/mYg9ElIgaZVImV
ewyEJ9kO8/MpZU2DDm8KI+mwoesRxF83/j/lHLr5ltCR4fu9nqR9/uu0h0CcdeFwKeFal1JV6ool
+W2RDe9fzojQKrog41uc4qcA/GIM4qGeMiEowm5mTHRle4DGCtqQpB0248HaZirJLLDzhTGiQq+d
9f71uv4rOzcRyH2csi+fqgEClB8sSj08dTvJFxfR1jj9OHDszv/y6F5En9sCkW58N+bFwlNLIAWJ
49MqX6FuwXUTyf15dI/pRyWaoOuMcpRoolsPNWsko7ya6xJsmvesO1dH4f0ISjgFZpRKa7aLsTGh
mcFoDY5Cik10OGTZnuvRtI2a4+wNPXVksiGINYt0n+1ZGeJnvvFrH0Nv+m1IPsmKOQ+KuRIr0ARx
Suhmz/tUOLwGMnq66ZliRFAXlCiL39palSUrJc2ioXn6qaxzQAPiFtol9A83LZVx4GHdAMZEcng4
EFdEZc1Wa6X3yfz4pZjXn143UeEUWr/i1oykF/AQE3WegCXDQoEgbtX3XkuCIQbJ0SGMjGgV9bZi
7dYqvRpXg2ZUIkOfqk2z6HXGWMvgn8SmT3KnhwmqnvTeSmhG+AzP/vnlLe3mopIdrMx1qaiDMPyO
rqPkWiml1eGXn/uOPb0xsG6sKyQaAtEwzTOl2aElBaet1bwxgIqr0Ya5gMgRy1YjWldjTJb1tCA8
z0OWPS2GWxtm2LRHyJwItbrce5ES6aqJNlW3NHcYa4Hg7Yq6f4Mi7E7iI4xTvUHjWyVB+rI531NZ
zsBuSlGRaSNWJpZH5XpOemr9myVOIQQVz/iczJQYbdUZNn807+qVzoqOpSn+7XuV5Jn3/CRlZ3n6
kxE/vLnMz299ILXCrAVpqAXcu4CUlblm5jpIfqggCRjXOOnhPu0WyPTE5x8ud33VFgxEm4x/oWuG
EZ3DRmFhLPTuU+hqvEBPIwJp9dmqCwadnxTTaXUGgP+1hFoJT5NFULPUGEKJuONDpjbQMfv/ARjL
qMeAKatAgaeCOc9RKBgngS6Jb97Hoc4yb1A8d+7qjb79iiO33czX6HqLNrosjqF9iia51zAHbv/t
awf6zuJTiiWgldKQhC5ApwNlOC86f9+vFWGBRPNyVir/i7FqI1TzT6c+pAq7eb3//6rJTujOHGVh
dXKyQAVVIZZZOIVI4TIJOwzgJ8ZP5gvQNoYvrCou42Ka239g268lrEY4m+GY58gQ4/B+rl3bSu5a
aAPEjSr2gAr0a8ysqK9NvgWp2jVeXUxtNWIpwLJxrt8N4O7iYvR00aKJu/QOl/VUN8DgNPIkKAjc
NJK548vhK8bIe9w+VHQ7uIiY9IdqKhoqR+vDVfDWI6ESFp36QaypabJMbvlruo8J5aIo0aBRqS56
MGYa4UJOfAUD0Ib0FXVCZJKKkYciJOO9a+fYmweyEIhEG1+E4+l55BvR0cnwANruQbE0jkx2+JIN
I9SY/XwKRzooRhsvDq6dwdM6VDFlcV21GI92lJ8G17o/V7CZRoBvJZ28Jf3LQ65f9AzHxLsW7Rag
e1x8iJ9esK8KMzi+RA6fqT+Dv5KyiJF9EfQbL4+B7JBGlDVGD/7G82nEpMGvNzcuQ1uReQ/VOO4s
stZBzN3LKaOqr7xlLB7BKxsUn3Y8kkKX3I74cDaZrkoEHIcDnCPpkZa4mHTvNyuM6lOv0y+LCNWb
5yK7mlw0JkTFh0RSsEiTRaUC5cqMIcSNpK5oxhd56XtPrczltwmDIruyZa8T3PRyDgu+Rl6FnPKQ
F4meDLja6SlKLFTaulblFR0oyTa6iu6frMSb7njJpKM9Zj37J3dMiRdoNJmryPEg+TeEsEkE2rvU
YM7a6lSd45FW7mGh6T1AAByuXBSasmYAQ0lxnhptbZ1HGY1+wDBzo0unkTMDJ8oOKHJkz96jaipG
H31oFnyFOlXa3qYF3GATeHFfVW2vLy9NvIZG+imyc4Ew+PbpNGU2oeGUgUVa0I8nrkTwOmltSNv1
IS7dbm86mse+xAqO7BUaDzK0KvQDpBqMCoPgnDeFT5tzf3sfuSjWTjEBYQuYxTcABGyGYOG/OpVf
HmanGCRfRLDwZn12PW1ft7GKy3JGMPDOeOg6uoShhtVKcFCu6FlSMZWHG3Wqv3K34Vn23DZEpmvg
3IphXs55Kgv4U2JJR4cVxZ2xoxiS1iquWqbB0jxdkRF12lAYz3HJHZYcglyrEeafHJPi3qbToDwO
qGx3GiAEpL7txuCGhIIxca/vlsIsYkRzYa4F2jDTnhh0SRObnxagERHsZHlHNk2STHJEMHVPid+x
U9DRN8udxx07BUZSTIZKamS7owPfyaJVcBH4821AvZ1i2TczjSZwjqqUH2K2MhUu9ccST9Erw1eo
8lVuQX7N+nxcYd3xMKjeFl4DHnG8mEIxas6oR59nYJ9MrNTK2piJlJoM/dgbw0gme+DC228T5GzR
li48KL5eLMnJ7gGtGKCpNI1g75opfolh7FVJTr4ezMHiFlnge74PpBNa11ZO1qBW/5mTY1ewlk/7
8Ko2RSOl2pzvyy1GLkaUFEu9KJct0zHT/cNIM5rFP2aci8+HBUffKDWlnul8Etz+JXaUbPGjDh33
sr9Edj1rduDXgdNNIanMyX90I7mkxNBuHfZwt8itGIgaNAUmxJ5TSD6t0y5HF1hRmZBUbgmpZKnb
4fucORrCxPMGlAetyu+8H1RWmst5jQlGJsHMIAUexYhEPb26O3PqtL0Dzq+tFvrlUvWYSMlWMsOj
QpIGDB0L+4lFj4JWS1Mngaf5LIKYYJ/kTTxkgZ0NkEhLhQNfXIvA/aaYE+P2yt9mc31vLhxlx7KE
VCXbU0aZXiSiosll+J7spFVK0y/qIjE1ka9KGXLx+ZSjWVSfNWDcIj1D9uEpt4Lsky3NJTnpCoMC
yY6FDA+tPO7Ps+QTG2xSXsFYiWvk6GLqUfSls2I0UFyvt1+Czxnr2C5BJ9reUw5rVYwQIVnYdyCR
4pULFGCUjRazc/J5Fy9rcShID5RtiHAsM3CCd6TPBRjHJh7vqUs6BGDX/MeNTaYCq2GgsEF9B/cO
NwQyxzWczLk0/XReapkm9SmD/ZJ5xT5YK1HGk9iL/AoHJhdGoBqrvndl8GbU+Xn6eKzJ9RBwvTks
G6elnljH+a4GTVMNHEvuNloTLb8jvgalS8wuOtyVpWa8Hd5e7YRoW0JEQxIECqVtxeGPr0tM77Ek
3gEwZ849j4BtmNZrCQYRIGtUvSLdpvW9nEZevgJwn5YCmIMaBUpsTXqSv9CzCtRTQQpvfqNwh6f6
BXSe74L+9qW/UNlwqpcu8+dTbEg+Q/ndFpjijSBAN2uEUOLJLn6UZMSpKGqoCtVzabLczS5Rgmwe
3Z2T2YNxkmbSa6npweMkN39xzTepEMFIRJH8Ynp/gTtmwLqtg6iitO1JpfYLEQzWyulTQOqp135F
KVhWJB0pN9mtmwtwbx3jJ/3wO/KnPqC9EO7lJR7UTiJsu5ThrRMVZogqC/qtdPgvpC/NuHaZOZFK
E0MxHycIpI8bun4v+eMpowzdPvskz0bIpFt1X+yAM/oBtVeC26ZyEcnuhj9xYFxXFO91XFqaVyLO
GzkTsiz83kdDxWBKnyBuI23hTJxnCLZ1xv26NTHIygwti8e642iC8taBPuKnNBkEapium0eTFQ5f
8A4fsSN8k3I9hb9/3GZ+RXYmBpE3OCapPlFsAal/kypWYQdBItZEmSnjebp+XxjpAgc0m1A/WQ62
T/Vh98KeesuKB4vFyrvLzYEuCfpVUtC2OcokHgpuRqqajLrFM/J/SZUSGA0G82i1e0O9mUkItyCq
le789PlxziFeKNfWyrOGzqBAGTWcfHvBuwMgunIjX9nC0NpOcnT2gRSFKGLSet7fDNulpW0lz877
k+fH56FYLVnXi3AlWYqCPvyRNd3V3tlnyf54CGFgeBMAfnqDIyth8a6LYZUlHvHei1Ynm/SGexQ4
2Mt++SyDo0nWDEqSRuUmbCpHZvcnbepS37E5d3+opE7AYW8+wWbZDEWvYPTLHJubM9TVJnbJDC1I
bgfZAB55esmWZUdLq7WsQkIRxzdf+4JSjLAXR/BtfFHHUFpM93rhTdVgG/+HoEULJrYreWM3ME8k
oS3xK7kMfx6o7e+S4LujgLrJqCRaRp6Ccf0ueotgNFdFVr1AGdqcivW0A429evS3n8JMbKQXaqw/
uEG8d1FaNiFvp+VzN8U++dModmgRPmloaoAUXFyLMB+Ich3cMUrljLOb5RB4AakigDG/pjRHy0Sq
/uUAnLs8TKUuMDWeaZ12ZvBOOS1Nj3fUYX4pVUhB4eGC3u38DrHt7TOl+JTrJVogz3tzQpDUmtZe
tW2RWNPNX5g7vrXirTCnuie11eY8py1drrJWY/ClC+/QzMDGyUisrneJ30P4x0AZc56OFHbRRsZD
zJjfAtyybIUwE07LKugd9BRqi2nU56pSyvlXQt3pizKzDnqvSYy2kXcGDXpfRrtD9hktW0SZ5AL8
Nx1yWHL1hEaTKKtzl3NSmSR0MrhMadyQ53yQxsM88qStiDfseCMK64qKJomW9ScsJa8FhFKI7xLq
Cg/erCd9phkw22PvA3HZHEqivOrNEorUsYC5E7x8+2rPvRMaUv9XtCJNihGNQtCavNRgu6FzbHyS
OfhCzuQ2igy+VuVIHI+Z4wB2UZieupK73GSDRrYkw6WeFvVj9nPhl+m/MWPFRUiDmG4yZ6Bwz62X
J3PXbml0GbCRpCFTP6A4KIgEyXVBaNL5zBhSmSOlhO5UkShQn4nvlryz3kSxtcTP+4VwO+CU6QW+
gOmJh6XY5bYQgxYDdL0P3eX4+FwLqzAy9BD1tJDXio3icMWmlaAX3wfd94MF2codx8zO2xYLN/62
fRAP0qdg6PNRcRESiwLHwtpYn1Od83cDFC8+ycvX46l/UNVZzl0dRSJtMpEsjJlKwU2m9BncxhHL
lg8SSXzL7m5sJLoFi3SJh5zbhQDbanIAeBWkQIJc2r4mJeewxiNEuH0zRFa5pFs9DfVak4KW+ctj
r589kWhRKQ/KN6/FhyX99a/7UJAdFYS4SyM5ZDlP4AE8ZK2qWhSdbHfVEhpDIYwd1st7RFn4hJNW
bjTWMG3EewBhjHtmshckzZdKFCGRNtve1reEVeyCgSNj9NImOZ9i1MhjjisILvz2oEPV4I8CvO7S
jm9JHr4BRHqBi/r9DxQggESTLVnZby8wZcB6JEQQXr3edEJHHom1iCGkOdyXt/AgUsStj4RDsM0X
S6Tn3O7/FygHVnPZ2jAdsP3eyMEgZZHak97ArU7mQyjxjMavPtFkkrsbkyLRYK7/aZktzn0ihheJ
oIKbhinAzjZA3nXkGgIB/xXHtipVO0ferZwVOU4PtHk2BYFz8Bz5EqovAGc6GYxufgAcVqwYKTe9
ld3oAlugkckDlCJifS9/Q3NCDkJDSPQ69P0u39jNZdzVnOfYt0JvHuTDFZXBbPBqCWUmJSyS0Dxw
QeNKFt7nkxh8HW4rT2VbZgA4btp8kqdgZSCbqoUdaWwaMeK7HVTadPLOlGaEAuVMockxVR41qJOx
xEkz1uJRjaefuMQfOiAk9Xw9pvfhJVkgq76jNmgqvJFOtFNfxfOalfi6mJV22m7YbqSXWE1ooNq3
Dy+kJAhJHeDtcNNasR6N/+ntyfObO67yFQw4uHjXRCTnZVFCuartvcxF8/smNw3ApJ8mLyy+CXr1
fMuyuPFxilBPsXzztNIaPrrn0qE6V6I/mGt5MC5sJz8/63A/a9nvkpXTW4NxhGfqR1MSIM5g2y/P
d1LGHr/NXOMdrKHURm64T04Hc2aoBJC0ArfFMaNrQUOR96QfzIsuiuxMcv7+6snSk+yB148uv73d
wBbm0L7ybV5aUTL+jPUiRuUsDyteFam7YaSy5Kvz7Z0zYG1oawadV+NOw146q6AWimo+wiHDQq2B
0OfsNm0rOEXAOp+/E3ZRArn3Aru2vimm+lLLev7fPV7mJYl3+BnMHHurHfApT8piztgF+li7e3b5
5rTX2Z8eaEYUJ0rO+Bpqd0SBYIwN18UBVrEM5AqN1hgNCaT8ghtd7wne2+AYTG9hYmqkTeuvHJMd
rviRz/XpEBUpGulcqqlt9JbyWQo6GqKLv8JTtMMz3njzroBtRWSZmmXD/UWxqBvvdjRielombjjM
ogI4SYg4e4e7wwDeTDIVT3Ebx22KnuWY2tv3zRO1pJ6cesA6UWPrUPOm8RycLMEkvjAb7L0yT7HP
8PDDf97bQXe/+uwjnX6TNoo30Ti/7Ntk2sqJxiHccL2iwmOMyA/zFeZ2mrqE4e7LGQJbwUvvZJoL
VWpXzFwW9MuQM3vpPTAhQAKeyZXf3syc9O64MRcVL/nokDHxxy0gYwd2rWI9geTDR+ZLojIh16nf
UP+uwgAlWXkWZSk7xWJTsLKL2yYgZbw3NJ0f+aFAPGvYji1g9rqU2zkZQqz6RsT8rAzbpQTDEY6Z
RGRu4vafpyT2q69Ez8wS0yVVMgn8cSNiWeJK0Z2qQ242iJh5BJhODGZCdZkNAU6wPyTz5zXNZVUn
FnQ3yiGPWeBY6fqbcBAKPT8R8MtiWKEYas/NwQqKceMra59d4C7amdydG4s9rainIlim3IQ1n6t3
+Xrn+Ii7aWIytY8UpaOYaeT9AbIMNcWkfASrrgBNPJMGw1zgMq58mwxvRot4JhFCYTGMYVijzUri
nLq9p0sYQ5zmrLgpZd/k+zjvAxAvVQfVYRsfu6h511us+J1RAXbqmWhy2sUqnCUlS+EzAIGxU4Bq
Pp7NKdPrBsP0EVxw9aoA+6NUouz9rvktnitqGzOhMU6/zcWWAXTG+QZlChbeGTmcjsP+K5hFs9yz
t4CuRMhbIqMmw7gAklxvMMdn/AHizZtDdwba00ryxoLojprVaPYd9H7FNoEiw36acjoGbzuU2UQ1
PPgn6A6wPjxjvpIWI3CyZDaOHbqOUinTh7M4QIFKD57SIDYlvMHo/hFxsjS0JXI9ryjbvSvZ16w+
Teg9IiJ2ZQdvdPRT7vY15+KsHihCsMDHNmZln6Ctbw0v//wkuHXbpNciKmJ0PcADGCaOZJX6RmT1
Bn8IOCg47SDkti/JuZ6Mr/CmRcp/8aHO5YJICU+zTBLD4PWdoihC17hh/ZVots4Px533Oba2JmHU
dWVRf2tvJoc/4RCKDAOqrvyXAy0BVjLSFU2CfQLavH1q6D+lW8Ef0vDmrvgrImjl5uhc2N5Dx537
Oq2smrN9rBC5FPCUsudlwyQhACg0no+kYZ5PIqHVfnmAOVdfxMTI7t/4y5ETY98vxXBeXNnKLNtt
7ovwTCQb/Ivk/r52ontlUrAHoCFn2tHn+ui44uuIbyD6xBGYYSfheIndCR9mQ+UjKas78v22guxH
vrbgiG1DEWjx3RMcz+MjC/Z5W+URndHfqu4GSlT6h5djuPclP3495L9A0dOgY2+3kfALkH1ZVrx/
PwfbtNa597TlNj4rEjLHitD6M4mLydeNqRuxrXZutZzVgbnaYJwx6BoBcK/gFbF2eA20rXbrKj+m
LC+bz+GF4ZgadruDG03qsza2vwG2l2Gk5dOjMy/4oEwFfMujVKzA7EdCIjzgq7FjYm8oURVs2tDQ
69Q1WCRuIzm4UD5G+MFDUIZb07VA8LlOeMEvHf3v93quOpv1vG8aNpQXoaN1PVgyEDCEKLMjJPmJ
cgibincUOeaOb/qQUPSBGpMnwp2CQGimL8XkcyqZxDXEzE1PjzVncLSZfG4FjmiI1mtEpNsEI7/w
VZ01M2No8+TdXyctNhN6DCJ7qa8XRoRHk5JCX3UlkVLIB4gDCkeGT/KV2XdypszTdZqi8ROhD5iV
/mjjoT1ORtfADQ1yZt0ljFP7+IXEbfDlfh0U4G6Gd1d95s2CQwjw1CtQB6NAjalZPGyZ2RXoakO4
OvynXqNzl/dvKACEaUXJBVNQkjkAYdU8XGFzIbgWAi3Mrgz7bx5AuNjH/HOPe6f1ppEjH52zLrWh
NRLI0Fl1vnj11D8EeZCPnja1EZZkrlwFZfX+KsXY5J5kqvMILTqVW23oxByppz268VoJU0Tm7edR
VO8FBTO2JPsDt9+/SGuVed5ss6CUJFKmM6rKvfQxDcEivABrhTZkR480H4QFHLc2CcR0F3VHZjVp
DvpOa1fjd7htbr+MGwatGS2op/uFDp3t88FYIyNxnVeeS9NMzhuMyVpVZIcWO/ygY8rkxFno+kVb
HLRWjStkMvc7NoJ1DrPZPEurnjvRoFblpKdXnGrLyxpR9S7vYQ8HIXblo9rjfpBgT5RDVTkwLq9W
HD5v0+25/c5AXrGPGVVpWXRWvfl6+2eZFlLPBkvjZZ32VIZoy+mz6Vp/pvcw71artHziAXzAFUgg
AKveTK3DHVbXe9NfummXFGQRwQkXPXVjSR4RX/mFpcMC4D+6j2DJw4D67EAkX9QxXaML/MqvSoAi
RH7TI/ksTU01kOWo6E9SXSvHpi/5ke5521vpnJ7jo58rhrpx+/pThvaBPJ49VmwQTeHgCqhbxapT
wFeoAYB9dfaoTH5j41wMLB9c5c56oJWoBIAWLwwhY8E8u96gE7morz9opqj3NW6ZyMXEmekSIwEl
yI44ah9yN9zidiP55ynwxS1MampP0eUhkHEDlhxg6o2iYmiO0jgLuyG8YwpbpKygBKUZrp/+vkh6
NpdWwy7uhA3uWw5YFmsb69qbCt5e0urWafMZLXkqZUXmIkLkoxgyIMIhWV1M95lz75Su1uJ1vDa+
/hrAHxt1tN33p7HQe55S2r9CfhEDwdy0gXjuhUg0DwVkOz3Ihp3K97QxKfyNIkbWEpvHL15r5cZW
neVS6RTJbs7LhVh+ty2r30EQHbMLvgi8Fw9IIDYDs68JBfgcbk6/1/9InzNjSN2s1RZOVL5AIq4P
29LOpiCRJlOMh177KqoN9x6og2qa8rVfAYA3bpBxMgHkFeCq+huVqLtLh59SrymngVPVh4MG/6Zs
tVm6cEzdtBH6rsMlH9LzWNwxt/pavqW+U1D9GITSFgECy2GW2Dsin16aM7XjeBqJERB4i0wlpJ6F
C0Kyx5/xu4Usdb8w/XxcTMc2dpIQu4Bye4lsHjHiGRf6Q0X0dBzwVpLxzethuyfZCMScO8jik0ej
zZgx/M5L3zLwLKJfglD6A2V1WeqCC0MusSb4/iRXvE4SeStHnj325GEAto0ep0uQ3ZfZRrmdR+qN
ER1OMJRj0y+us+vN9ZDLB12OnzQfx/YGAI/ISYVYXL2hIxgHU6zuBIZqsXuzrdPJacPTwBwR3kXO
VqVAbxXROBvGcAjFXMqwZ9MS8kqRM7lox0sbz6/p0iOrlBICDpRAStBj/Ct9fA9GrEA8J6yBg4qy
PuzPSX0EgeLwX1xlS1Owor71YsOKRaI6DMQBEFtnWhvios0eX3ou/lhXEygiN5UAxHVtvrDOOmEx
K2Mr0dXyio9Ck0qSsQsKxLhs5d7awcOZhjgYoHiiiBVgzbXH41alYPziuNt+HpZlQlpndaiyeHyg
hrJSX6kU6JOKnK7HBSbMEmeOhYLr7wB9d7Dyrg1vRckGLZZY6p3zN8CVhYgWaVtXx/S5Ggr4j2xu
GMF2Bo9LjJZMn3MzKP7OezuZrBGIy2sOCzE9C6hfe2UHS/bh0ouLQcNHfYO9FFRnLY7mMhtyqSGJ
retLft4RFY/0unMUA66KQcywXSwZDD56ffE/oK6wjoFQx42GV1eTSfaKHPQYSXKh8ny89yV7NbVr
c1y27DlUwnKLjAcmMtLYWheEbWHcTYl5y7j8d+WH+P42eiR5bTyHSlypDb5npao8LFZCeH26Qft5
wydwCBaSbXYfS7g0Yan7WWdmcmYEFXJozHyWTua3A6Kwh32Gu9uhzCEkDx2BM+OuvoJg9JuN2qnF
B5zo9xbXXmEiko9nCrd0BrPmNqBibpK/PcYWok+lIwee3gbAMaHgziqnCacGgqwLpxAnJRy4Zeaz
SXa++bwclbhBseGTwQcAKfsb3peKInVQpuArPe5OdYvZ5AXKqvNtz1vlnuC/JX9LDcgCekYMKXKJ
v8Bw8XWHATwRrgf8akcZ5KSkeraXlRC0iSc6PDrUsFiPSroIdhKuIfj0ktEKltDyZUwaTodvKjuf
mQmIraYB75OdaFzxbuV8wwXsHeVxVc8GjF6X4gQPoLLyr3qXD8pRP7Dzs68JgJB6aFjt3Iuj2LY6
BYMEGiG6QYi6peyjghCFO0/8QQzuo/zzxcQRWvhat2jqhWfXa76wG4OltgQJprVR85YFp0DUVXKo
15pOku9RxEOh9rS6vuEE6CgoNIaTaUuiOSzLi4VglSU7NHW1543p8btmxoe3rRkO++B5XKtUYNGO
nLKvBnoK4I0uFmWW+BTi5nhPjdvBvZJxNFzfph1MJ80BQsAj9dezFH2Uj+y5wZf6f3RYB28yrGvL
2+PgbQ561Tyr7/J9VGrPLZZ7Sns9LThR7IUaxndUh4kWSpkxlK66yGU0OEtzFGkpecllKB9b4+Hz
29Vs2ZSH2un/8brGNsBLMyqGorLNTljGqtFaHnJTfV5TlcXANnO7UH2prPH3VZTUTszNNSCf9pGw
3cDSWZDO3cPI5nDvqUZSPb52cAAHKFt0FhOJ/tPWRQ7cX9cUfHbc5f9AsQ2C6r471gUu2f9YA45B
ZWpvshhDZv4sUwPoUlEOcLS3iniAoSBEXly/XCoP5cwN3DK6Gr7TMBEJh9LYlpAutzvKwDu8EhLf
DbOW0VKHZJf9RoD81TSc3j0TAVo4P+F12/un2KcrvvXGgMrC4mTGVeUowEfIP6ah5pYMGjKf9PSY
rcw6h8JxLQ6Jbxex/x/EK+/8SutwvoaQ+Vsx+28IlrcrZItygX7BIgmR+xuhXUwlP0SuD0UVPab6
8VcUJJBOYhMg1v5pNulgZh1RqyaEOO4WlRfPzpHekvPZnC1owkuG8O6RJeJuTqyOnmp2KmHu2DzO
RHP1NR00QvOF8h0epYlDKF6i8Up8mTekKcd0sod7OSf7eQ5ifo3mus6Q85NXI5nz1iFD6cM39tAz
O9AiPDgRZCAlqxSNg+4nqp86mhihgE3HBhGx907uH0B0aDB2F5Xh5zIIHuBkqfpLvgJAVFFqqywb
c65NV1+XJZl2nNTbUXfOqtZ0ktyrwZZDXSBiUs0rKBPjGhW6NRXoepVzi+nHHkE/xDGkc10aogje
f6XqQD9NG3/uh90XmNeqe47ow0dvGU7RBOAc2A++3WuPr6KT4WNlY+zoI5dYJ6SLsl7mosdDNOkh
+jEm9UrwyhK6ZDABOE/QWA4sY33kB34sTAzoW5iH8KthhGqM4M/ZDseD28kmnRXv/X9MDebYkCp+
mrLQNozZFI2sDC9hDw+5qVFVTm+WTCWgRm5frvyyPBuxwOoJi0G8TyNFfZY/mb2Z7vQcQEgROYwF
kDNZRF7jU8eGZTTTpr1cRx5vopHVmLPe2LtZJHtEcqITv11YgLG0F6JuLnU2fgOazWnmnQutbdGD
1SCuKRFqy4y5JNyE7Rfbh8bXEFRWxwIyVraxoSpoWPmBK3aqY/l1nSW+VVElIZLmdRwMKkuXUqgI
c2EWmmRrI5pBGy09Ki7oLf+GMkRcg9QngUVFOufg4JuNso2TXTHMijDpkeMr3bOM0zeIsGXTtCR1
DsCC+MP22HJn1NbfGv22XPz3SQZHrxry3XwE1AZ595W0wKXHm/BUPuk5k+Zx5+JFpJAQHGJdew+G
UZ3koe3URSMsojR+gVFrgcAUXGULWg8jgqTHdLdbmas9r/ya/yJUP/UKwaw4CFLNKcRZwEdiqDvK
YzuloyLIxEGEwSYUZh8I6W0LtSSNivqWsy5S8otyJIaKRRnvccAL4E6nOJGFZppDq0M6C0hn1goA
NTsl3SVYt+JT9zHZydbFIIJTVM2XAcgCMWk8CN6nW1zlcRLMwdHkI8WVF51NayqmImYWc2xJxxB6
Nvyv6TuFbTA3UbJlwbN6j1HhF9elgQ5IlkdXTcXo8bk2tpuj4ZalIAWlf2g/Nmv2vK1NuePwaE7I
hDQH+DSRNN5NoT/TwZgJpBFedwwA5hkSVVq7yQ2qPg+MRum0rq8B6FgPwnLeqRWoAa2j6heQJLdI
RebEhXEIf9yKCuHb6nz9qnV7Tf6gSRzFnb0EYR70xxlwRNZJwGBsFxXIO7zpSH0pZxaOzBbWH7Fc
Pc3kyPAaqAeEiNMKUr/j/0hUaJ42J35yFC1qNPMtfcWbewryyOSTJAW/cAv+OGkSThjZJRRmjrCy
z7dvKnzzWSstNrIYKaP8ZQGEjcDu5KsxzkaioetewLW3wEOC3HVAd18OzUw9J+CxtNdHTu3B1n/I
GrZcGg2R/hqOqeUh5l3R9Op0KhZ0b2yNuu9whs7KajkHbpbFKOzb+ye6d1hrBvO/TnOweTJ3EHdg
nLpD6jTYELJsmgk6+ssSBWchDiiTAdjWlMQ0t2DQJhmJGcaRgg+szy6fTSbEW5m3C5vGStHViN0R
JlAHXgYjDvhSsaCYaGkeAQJFYNxOs1z113bI8Is4VtM7tOyZf3ISrcHs0JefWIONHaX9TApj3+4W
9AFAGeGkpQaTXI34ZIm/Gom7THVezVU37Ejofywq+28xy4xyJvoq46x5od+n1hKRNZYGm9DvPTLY
qQhn9aFbZVIr5MIrH2LFRYSc8aM/fOIITg6Z8tryxdZi+6rlKgkf2xcU3XIPFJwpbIn+TqgQQp0c
czvpnM0toS+ro1O5soiG/2+5vm5H7wZk6+eC5KR7/qyWtbKWcfOGegi3gBIrMDDG7NIi3H3GSLFU
uXQFuW8TEmc1IYsGxj+dQDxGwLS94m8fSr6F7ZzV/Q59F3fY6T4eqEllr23xuVEX1WY3Djm/nhjn
3+T0tJqOqjCBnaX6G/4Nmdxb0hPB7CDYbzFjaWn7FCfYFji6OiP8O21DQr2F2aKtPWQBrazsZsuK
ap1FyK3h98a9evatS+AGTrdrEdSbXkZlB6lUBcx2ZU/FyIo9XPotNCBE9xSIVpzIlJ/5Zfx8nq4E
evi6YTg4x59EWj7LZAtDt90XgtnBJ/NUEO+kG7stzg6LE8TZtxuoEU3GETd0OOHtPViNm0thwQq6
/HR34R16C5o7luUSSyP6L40oJv/gLblaVhBmTHgJVCfLZMpnhNfggoGduT9hS4nz8Nnc7vJLqIOs
SPRYQQaoem7umno1ETl+jeO2NInTDRc+tcfntMKhxHF9jQWKOxsO3eYokRqice4Iqdn8jXDjMXn0
+8Gyn7qjRrsckHT2Nb3njMpz9SStRMmOFCyoSKr9Lb5vBWa9OBvZr3gM++pcIVai4gsZMShe1W+2
rkaVOs6kdVOfxrVAMawBouxgVF7Lwi/W+S6pgmfvODB5qpljp2H5vNyLdojVYc2VV/d+ppFKaHT0
9ROri/8iqOaXwEwT1USnPloVB9Vh6Fgr30M7V6dQvdZpE7HuiQapimqOdQTDeFbhgTl748m78TrN
VThd0GM7e+Qak/hl6NxkhtLUw5KEoY19erESPHO8YHmJdTvWQq0xnjR6ZJuxgelaqYPztQ5lB2HY
QJX+JTAdCooDXmIz+MtEVSf9gfm88VcqC575lbePr7z90EOjfBlVF5nnwRHFa0l7EMvGUKOHswHI
yVtc9s4UbgEwSyfD3SkFqP+dHIqeMcydUHHIgGWWvb1fRlgh7b24/Q2DybiTNp0PoqqKBju4QpDH
xgpPGKnq0R/VCvjspBA9sefI3Bb0VNvr9f4LReifIZtDPUVmAryKyK3ym+nz79IW5dJD0G/zrGTA
urbGrAXEMe98Aod8UU1JEY92P5x2K05I70SMXufCRbXW0cOoW0DTuZ2T8b5Nk0Ox4kpn4iWYhKw/
nlYHqnJWmLdrZn1DCfTjMA7esfc/BVMAbvK6YBtHQKRz/JqyOVp+5f7CNz26APba9opgPXIdN3Dt
gTjEklsUq+u953fz+Q7Dt8veULfLvEg9CbkHddLrFqH3toUgT1zLTgDYN8l7zwSVEFnslcppXeV6
fu/yk7nlexLQTZ7+tHEvucFIVqBWM9W3GoRZq/BtVqsJpv9ZoLrLqKIQTocotw4Az47vpMAEWdV6
VsDTAIFLPI0zT0O2L4HB/8a78xjmCESggyy5GnnCpyA1vnJUEyOeV7JDC/QaN/13RRhnhP99Fm/I
NMl70gsoR5VAy+XY+oUh6F/TYnAQN6Az/WqxmXdM2ktHrpSeMxz3XpaIVO5dYoTq08uYaMbuzjEI
xmBQ0vQvssKez4K0efdjG9p2coJugI7cboy1INPE2YBQB+qEZGgV6x1fWYBwKEyUN+/eJFcOBdtd
qztcgCgpE0pNfkN9Vscpfvw1r4DJjaX96XVpmaMSTykj3eziLjy3w3Ca40JQlhs9RY7Oq7FsmbSM
K0LVHciglZHt5syh6ao4FL7xqTR2E6Xf755VlT9aBcp/vgVeKbwpJi7IH92BbPCDDMHssRx4UUlY
YmklWjcnYaVFuvmVQPevASC7ppSpHNde9Hkww4cH0zwUe+7kuxGfJajMHLtNjXkNGJuUFtWSw1MS
oJXpXSyF4qpIFuiFU1EkMOoXLA1xRdEG/Wkp8bOIQM60tcwMu7LlNc8Sm4v4mhtWxe9sZoahrB/h
IN67RchIwifvEkt4oc6th0k5nFoIhhS3ST9DqUBd4VDnf4iquLxwA+KuCuS/60aj4J5GIRPngOcR
yLukfLS4OF4zVb8CSrqLqsv0P1W90I0SEkhbagcwclGY3/rYzhCIXiNXikUVKoKC0G/99jO/J+M9
/yz0yZOLkHBjtIUZBgHfKK8pSWqMmG7Na+AC+DFT3j7GjTrWIfg6HDZbXY6xWGKGr/oWdsOhV+rV
UExHb9+RZN5x5vBgmokwQtincrTrVJ6CZIyGvEGwJtPW6iCbuDdMYlB5KcUscbNvS2uriTniB0Bl
cJgCDpw9BkOqIsl307ZzuoRlCeYQWLpTwVsC9YhBiPjWNi/IRk9Rhdh4Wpy3C4MayHWF12KfXRwa
A4q0wwPp1KKRJpa+HKmRS0fluUt/00irL6OZLqSaDCUCmnPzWzBWtNiNqmsTqtXSvNZGgzrvtKYf
dhol5MPjiy+EHADVmC8yJKYoxsI9zHmShHDtmmbxX80lgQ7Xnp6ew2VN7yCGJlWk0A04Crr+mtOl
zDVXMD92t//LpNFX1zLoao0mkLURh310HV1Z/cvVGemCkg0jVKPMXjxuNaMEF1yTf9WkwLsXznLN
b7puBdU5bHM8rPyGmIHYgWIfJjBZAmp2EomK4j6tKrtEXQ1U2e8dF/HM/chNspKDH8uQsBxlRlQA
tI7YEQP9CU2c6lLRY5GjLAP77J87PPMclySFSg9qkVGZgtT8H4qD8JLgIhmI4jrgTfoH8/MDZVYd
hDzR6CZ2F7vZAE9+mYx8k6lWms0cjZcGc2AMJ/Z3z0LLjOJDDvsQl33LtwltSJn4qtu4kNE49Xsg
+Pnd+pWR4t9haZFy3ZNy6eTvCdw8SkIXxWPive/+3vNr5N6WgCO7KcQNTcOYAusWLaOqFW6Sw3ei
L1dWiWhiUz8HK1zLVkJKEYflOdlHpzorL91TNG67OpMuLqg7lzPJlrFi6hj0jjA+9e8yFRyvKjYd
m279DIxmZF4vgEhV/v/kF74B2D7nqlAyw1Z9dgx358RHHqJPWlBJ7mz0a6OvpT+SuME0U7sYlEbz
TsmNYVddNqNxaF2DFC+PpwgnkT/jc5Mu2i5KVyoBgiHdl/mFeUMXxDvQhBqJde0UFt3ham+pCqqj
dGwB8UDOrWSO6TZGnsWGOzgiDIgbTo1imOoLSu77ZSc+d+n9E5U8OLye0m02FDxU4OARjP5VGDhb
0ykNdSMenuwRexQT8mskUZ/lBlb7b8BSt6CtWZqZ+eaBXVhLMppV52ekMVTurjMdPhcnAgyCA9Cn
muDtOgf4SqaVDb4rav5OiIIbezq63mID6qnHK+IKqaKrjEA+rBLlqvOMoy+S0BFpBmrm+SUD295+
/vH/dGsponTLsYgZsYXX/3TuxE29CMhNFy59ylXCtTSg2+UaiBDCdcizzPoVK9LKknnAOu0aD2vo
iMUX76q43a9FIy+KuE58mAMT4v9Ya/PSCqVA4mpbNlfSRcF4k3JVzr+AiWG7//lmeg4vP4xP8dfQ
zjJzqFK1X06PJoojp/MUm7d031Yg6Bb0WTEStD1PFqFKRgnUc8MNU2KB9u6Op9EHr7PhOjpWqlgj
fY+KQSVvpuliDIutSvxb0sSsgGHabIFfv8/LrKv9vunNn1+28jWJ/0VrHt74lLmC1LN2Bi1CB5lA
fxtaAiO4gM/6EfKTnrzBpJec3YATlk12RuCjz7brsglD0tAuW8QipHr2i3tDo9W4vWYuGXoK9r05
wTaQ1xEcGo7q7FJU2yjAstDaV3UHORUfpEJnWbpqCT0A9x15bPBXgjmzid0QitjJ7Ar45Lj3qNsU
ttijN0aiyYKQ3lvLHtwymqOFeo6I44C6DLVudUgYINOInr7n8w0pTWFpxASVRO7IfVyiBSwRuGEV
P1GVM/kYuha9iKBAnwDJW2QG4jB9Yvl6fxSi7A25jf/naCHaUpcloXnptrbdQT5D1P6m38LoeyEY
VFiAUH+0ubRsO40oDu7shQw3QDBaHcYFY5Ik5w2YYWL9E+xrHPwMVEMCT68D87Ar7wIZfbrXPq+l
nIF3ufzwmEpzqBySBYK4RSpAbMs34A8OERKIBOaDSG8DpiQBUuIR0H/ECGv42tV8EFEscgPTUTey
EYQOWOYiN6WG4U4buCiRjCh7hV8fdDSyeSQcK+l8Io1ZPuVh44MRLWGQsa9nAmOlbbU+FTVKDqiZ
xfxpwiz3P83uUROamhJnD9ZahUPFcFkOlJpDWNQxhigCcUk2D/9q2cjWy0NRK2yReCEhoD/kkB8C
6bZ842vJE5IJ3uLCp6qoNYCp9uQlFMYpnCe7YGBeqkOecSvACGde94Yr6WrOc2UyHQ6AL5aveT+/
tSx88IlRkLHx3w/JSxKVsMLoHCuD+8olHA91Rdp+cWN0UJ2TzezQ4LKJcA3RaWes5PTOGnQDfTsy
aNgZm8JgSrOuHgYdAIf5oCbe6hU++e4Wsn6nLipUAwu0RZrb+TMw7mYZTik6GyxAwheG8N8fp0AH
LzPkPhKNvJ6aA8dWjhyUSw9DOi4RdlN+/5rLsndXFQG2avpFZcO1wMvzGBn4em/FO80intYXj2oh
7nKRznfngEc94vH7/n8W0cu/3WC20RckPeHDlVdQLRxkr9ji3+vw4iuUqpd340LFakCxOFCeIFVB
yXfkudgJQJ6l+sc7dYdaPFtHZoh2hfGRkHSWly+fQA+H3kibLtAjoPg9ZnGLH4FdbioSFXURdfHf
CsVtnV6PKt2PmKQQ37pUd/NTgD8ZWKTD3y5aTYf1lSO2H7udrcCS2xpEie1x4Lp2h7KgYCOjOHcM
5Kq2TLc046h/HBVv8XBznfepO9q3rHQWVXh00QU2ccR+5yThT7p8SMaBKkXqxyQpXXcpkawKnNna
gy0TcJLNfSSKEVoHIktOVNQydcWa2uK/9rmku8MOEOAkuduyjKxkB+KmDyTMVi60TqWbnAINomWH
2bkQAXFEg9sPAhTUPZ4ilw2L/V7sOdgn516MPsRPUea/c2uyZ/5dwufsO/PdgijRFoMMHAKNIZUx
8qvvez1D5QSHIItbcQlNNYZoz+62+drjlcjWKwbtcZcp5oTyaiDcL+OhspTo1rTmVSjoa66CmiRV
cerrJE5N5SC/J6tZxdaJngca/g0LsTV3JNECpp2fXQR4C129+vkGk9tuJV5c8/KYhf13I/g9cxjT
Iwfj1UhEFInRxq532ltF2GTTc/VvVxZDZoeF8IJKvFJvgjyqJ6XyV9G8EX7Ng7OUEDOGTbmHIdeo
fr9pm22oF5nsu9xU8W3xAft+fXcTY8Hw/e+lc+cMUJdm1BiQh9SdRYo/MDaSy2OXnlBKrnRAt4K9
C9HJyI7TV9ioi8Nnblq8EJjzsZWi672SpHk9AQBoLkNiJpz4R7P4h8X5G9Gz02wfI970hVCWurf0
pUsRPkVLaDQiTIl74yq6yIcimo3FwFjbulgPbomOJkEWNheQlhaPrPCZvXN0e95ho1roETFdgg6V
j1klLJwo91He8idIN2Qhr791YaaGnstHBLK14MLqlUz3C4SJlziXcTzpGHB8tBIT6F55BASFS5TL
yAsdBPP0vxbuJ9pQ8frJaJQytge0aTqqjdusytBXhiADpZo/FK2E59ZFDNZFp3tmGW5AolAtzIRo
TSnaOGvoXH5NdVdVga9KdjyQdRbixDpdN3t+DT/Rk87ecbDQgw0oSGkhAp7m3119ifKFj2L2fD3U
nJIKiLlj9swpWmmfOwakp0u09RGf/q5pU/Q5dg1YsJxSjwxj9d9Z0nuSYARFR2hY7hT6pZCXFgj5
Z0GR598NM2qFYiM9tQ+n4xkUnhKT4SLG3zRNrRj0GT7n/fCpb7o5wDD76YseaXsXU1zDSQYtJnQF
o1Ltlqd5A8eocRpdopSLm755ZQQeTamMugG1op8LECiPjkHdry1LtVc7Vq+SOcp/e59udJ0RPsBz
tKD/B0lZBPLI34bqJTbJAH5s3iXcSC6X3aKvxiu0oGzCL/lNOpMVyGYXRpX7qRyXLLZK69BEy89a
2zY8nqWTlO1B24C5cs5ox417Irrh29cokd5IUUTfehQ3qjFu1Tdk4GOU+WQKgHdskiiG2vfVwREA
81pY+Bxyd2CQt3pwgkVPL2hKX/caZQkJO9NBY9Xg2yMxLnjnGRUcaACTFAoZOBjnCg3uoLL42Kvd
ZavAoqQ9KTfk99alOMcfop78XM3vyuJInBR+DddglP8GHwQ9B/7l1h2AGobVkNzCFcApxW66S2AO
qZi0JgQ3lODHs4yctMBERIEtTp21x22MTf+p3Lhm1/mzDysWC0s4AkbnIExH5X4I5zjYV9bb/UO9
kGRX+Xr8vdtfRpuB0j2NjZRahb7+JKsUJo06/2pJ+bdIF8hbRSLYpV84PIiaq+qlJuRGuKKg1stE
oD7jtZ8pOE0vxTMxIIIOnj2jVt01QP4klaVG4Wa+oxUblFR//T4KhNcv6nsVKBWiXAqUNoge/IRh
nc4PBeSMOFsBo/zPvborGB7W9mww4ErJheCBT7LuPNc/7uqbnuBKqr51IaUyQz0nfRM+eamMgtMH
MKdhj7JNcllFU84RIfgauBbhEZKSW1I/KAo4qnEbXt/q0sk0tMfnhebf/z4yGEDuXYcO25eRkbfE
8xDzME/CifYzN3C8WRi/VBBsiCz+9edarjgIlOCp2u+EC3LWWF04jthwUqKts653eyjB+AHIc0AM
kzk27SlLKJGQABTXnGRO+VSJNi8Yw1m9ftg5Z+rVbLbe+l/qBBDv1Ox9cG/loTVSmYeWqwvLlN0r
P9Gq17POc9FA7z5Ew3R/vbckJ+r92YcdxfHVcBHllpS0XqfHoidKDEMmfI0ilyZcWjyUdIderScy
YxG7vZ+4mJ0JoZ1t9l61oStcDC9QxxFE13FPXV1OmVgzHEGiGmV0DVpLhGjdJkXDfGBWdaToyvK/
oi2CPPXF+dUj4HDWcyfTXpBbXgrhYIJI5mkR9dGI6WQuQ9kOKgE8mIQGYeV0k5qsJurHFo+kZNFe
3uOpJrBGsdOSj86a9i2FKOb9SE2CUGaoN235D/l2MiTabDeBaVRZUxW0RR/frxvv6GSH1E9uDi7Q
tRTtdOqW1CBH0vW4SOrMBRHUaH+HBOM/e5r3HcXhdAct8mjtUwc5bYAqmC6rbWBtF3mPKymo+Wpm
BqbdpPUA53G6alXox8tRObWIiFVIix5QY0bE4wZIzhZGqvysvAMkOPgdtxoiHpVXAeAaexrseMRR
gPhH9Sm26U8N2hdnW/Rc+BrAW6YF0G2kSNYx8bRS1uouUTiCuKbhkOnwforytJfE75pfLGc7GDos
V72YZDmCzr24iJ/BuWBMJoZRS/6+oHTpdk+Ozmt8yVOPjeXXSYa11El/4Wc4oB4hw3c/6ZA1Mt80
yMuwtMSGGllJgVpBPBK9m6h2rcyltFXjVbwqsrYrkC1BaGQfEp8IL5J1BdnxmXywUAwJDjHPWfbz
Z/t6yZugtcI36HHhgL7A0MuT5du25JBLtIZyTydH7BE7CTp23E0zkddebWC247OG4nuSuEoEI2b/
TM4Ui2WGrDuykgUHuutcR6U4Fc4Q6lllk+T5pmIjCObWW5Mqqf9sm6cXsqQOwCiPkCcmdfBPj0yL
oonjpicMMqUG7iVkiuDAroxKF64iGkZtghwJ0D8b32V+xv/9i3GtAk/C3aiO7wVoea6AhB0H9V00
06zBqSynxUv3EMeHj587fjSdZMpa95ELmnHKTn3z8r2oCcF7KiLuovJgXCd7VIir9fJjCqBWTsxc
0wiVtM4tbYajXiXLTr9pygLn2kxEJ19HMhsbbnDXhVMYaE2P3OO9woWf6ZdT9+YHoxEnZ318AO1f
ONsLbU9UwMonbyBbY/rHZa66YvghYClCsixgwZCsL6QbsKEAF/072WtM9aKVIZEdKDnFRAkcnC+0
nLzLGGUi0leo9hL35QctHP8CXOJ1jQ1QiapyvZTmI72eVhxZm73P1MkchNpcSN1DxQ4edTH3G9if
OYwB4CETd7uUGt9eJyslqQ1eoMBuMrxDh9Wu8RFFxaF9m0cGucGN9F8FcZXV+MJfvhxj0IxSd9YK
xI+0GdhHJl2bXJVqShVb1lNemWgFpw3c2ZDG5X1wIwmA+LpkhY3/J3s5lt3pfXw5pNhbhewW5gVP
y+7pND6Y2gOoH+/iDs1rVe1ZYlL6V6mleqg2/v9uD/4W1lamySZS9UD96eD+uo/MjWEtfxbDtxu0
E14Qh/OL6w61y/civ2taJUBfAuCc/m1AcNMZ2oWVZg4dcrBsvMEP+VBk/lUhDWzibY4UtWZ7isRd
KT/HcEItXnb4DAtYvCOWivemQacsKMjcGy+u+R/KZrp/JIjKpBJmc17uv1/kG0f+pbFfoQ5op+VP
T9fWjsW7rCGh1NiaIQKMStjz5K89WzMiJQzrkxYePQUQOgwseNpDdOZdNFhB1nl4yTsYUS6EEs5V
HooBcX9ty67dxjy7MU2mXZ0D7UKgo1s7TjKffYPYxQUugOhdVXXP8R/uDpXnWLcT1n9Y1HboE5B9
/b8wzI24oAbDY3PGd+s7zS3eHWidGszuVrcMaSSA2ZA0FgkIbj4nT+S3/alRZwqKVo4ObW0O7ehg
XtR3vwCeaosR1nKPsy2uhusuOuepYreoiVhAwMVbCth3j985gSKiIreJZtwRhHUTGsxtEmhV12a2
zR51/1JpJbi1P1n2T96AMCSEcMRXhE46s7O6T6hk/383JMxF1eg8y9nlmyENSrk/9P+RCSlgP+Cs
eMfl5ycAP+dVKF4KvhEibhTBDvg2vQ3RIkNOhIf1Wa32/GJ1Iq1syTlLe7cT+2znLlEfCDXc7R6n
dgJtV4q3Bor9r2D+03ONasIxevQCh3lEaN4bhpIXdWTYbO8u/bSMj/FcJCUZch7lyrUgMnVoArG1
ZJAphSW15N7RP2mkXFmqtmhMbpOiiuTJnubtZUFOfdG78cHuXU1dNTIUXypxfk7eN60abIJJEqM7
xRELxeKUQynosnP0iOsQYJmcwVpRF4OcPX9KCkP/F9RebIf180IipiSFaFrSOeLKj2Fgn/IB8HeE
dONce5ZRUC+LQT2n73IB0w9DNbyEbFV2sEL7XKfyWFz8qI0kifanYWu6ba2gjVSejsZ0KXDKY0Ql
xzdUCN1Uc5qf3jYz4atxewATFVdwSimcAeGscqtwMiw+c9qo5ZfSZYpSrdlxI2lr28nlL22/2XNX
qjLAF7FUYCx4IPZxbthYlR24xzfj8/ivoX/7MDVgoFtDMnl6BUkRN7jVI36pJyQKrrUE5qLRGgo8
G5jUlUxYBh13xwZFvGUy3IgJ7xMjqet2AFSNJBiXWdGzCPHzee9agBhHBcy3HGeTYtEb5fjPEPVj
JwjL6WK2f+zTKyC+uw2r4Xq88HbMUiBad7NIzwT3MjNt7P4SxRHwUyEgSFRxMHAYkXMaqTKr/F2f
9ilNfSaxgH0B8Czx3sBFGrAgctbjqWZFv6Ds/8XVx+pFbZdnmLxxZmvWJwj2sy+HwsYNmx4DFJOO
FmQZKzq8i/yN9a8ZjdLoxNM7QtCDLn4LXFvFSUvti6nB/qNql9fWM5d/Nk1invQSVHpKQEBNcLOl
lfHrujbMiYmI2qootuW7oWgKs6uO8v49M8FP45WDNNiUuBxvndOYUUTJ1PN+ZY2G9GWl1YknHGWR
ZzHkNeYFVW/K1stisGYH75CiQpuKtqHnfmkazLiPOq1BgQDHebsWpeK8B7C6AlAYyfxNrRM8Zr8m
IK4VRbZDeHk08KS3ijZuS7vZBBlZKh9lNandyrn7LPe2lSe+TK8tFfi1OY11gZPIOxtpK194slSd
T0xAButy9esw9Dsq3gZPh3utMowUJ2PkFNz53JcFuuGb/4l/0ww0q42ib4WwfuJR+VaT4a8pPGkX
QpExbALwy7x5kCmQWGzAb8DxOLvgjwpTMglJtybC4jZce4gNQG1Nj/gKIf+32vbBYVF7dQ25qgGd
wcfSJFd9FaRxQrXq9muPDawLhNjESpyWJnzb4Nw2APiTl7NBpg20yY1ABa10uA5LWBvXAJu9gmG3
33AZoKUS6xwtYzrbbcrw2b0lqe3yZiPd+Vq3gCZrVdSCoJI4LZszivd/nwxvWc3vS7GMIRYXRSiN
90rEeghmknl1gFbgrqa9RLsAt0BIdlFUy26TEI4bta3Tbw0isAlUY+g880hpsDCibIEdL5nuh6Sh
RG/1Vuzy1nb0H22JNkmq8Zg0wLgRStTtiufHKEsdU8U+/84a8aZbIBHNoYbVNIL+yo34vDjxZYnJ
esOKYBH0h6eWqwOvkpE4E6vufhvdb6fC9HjFAv84349YkWP5qGoIU3g9AlnrEZx+PEuQxv387pN0
i9lZe1XYcPkaXsDTtjjIonp/dXawxSppFCDBoLwo9/SMkIw1Hnm1SdbGTlrhyUx1XQuE/qw7KzVu
qqpODY7slQkdd8cEEc3zDuq+DfFery1PgASqS7yDFZL137GtvulmPTdnlY/IXg/+IA3SSsD1ExAY
LYn5v3rxrNvi3hc8xO8mguUGnqbW3SAPJPUqbN53Kuq+sl4We9DIZgPCEUKqgWU9ovwpD9LIAuJY
6vzkwPgQ0HjHbNwi74Cse/WojByS3K5lJIXDqsCqhjsV2V7zpj8rS6tnTHNXG0a+Au8Fw1gYdDN6
BUjxt1v4+muiLlc7Vc57tJ4UxdAsWViHRVQXNofXKQcf2ZMxhHf13NNSGXiauR8iq/0akbo1e3Ej
0iZY16ycaTU5i47HzDIFkDcQwEBlugdPhI1868uxHGyXIukQ20XbDWS15CBqAX6+J0y9sjxlAoJH
w+T6BQMuaj7jlC/4Q5MN+u5jZIVbiMUGQ9OK6bfzRYHIabwYBCYqeMyFoaJy5SFVS+DRRAO1KGoc
U4kmZMqUvX/3990Y/8IygOzt92k4KMdZzrp1yTTWu3Iq2yCU4k2PzSFEhuxZaJeuFDQ4ckLU71fC
+QFuS8ax672z08mv8CUBjQXHSMeR53OYKw34Tub8Pg1JaY7+VSRsjU5fJy3wbTheJR4f0qTSr51+
D7NjDMhIJAtu0zIytYMmBezkP8odWgk2BojjdthfbhAYSDBr1Lxcqv3VoHGAevJU3KNUqwPOArAo
2/akoWjvmWITtFqPdpj1I2EB4K3b4Wj4yY14z90lvppSl1E2x3CFHEjIIlj5ImvXWvDGTIy4BYCD
WVxKq6YTRJAKaBsEpDv2lW61CckO+80yc/BNXZNlZLzVWUKj30q8tvlZP3WZtyNVRhD6+fjsMkF4
RegTOeIfwc9KxAkPVDN1GyUCWxt9lbJL8Ar2FNRCaKmSCI8pDSfYBWvypqpQjtr960+Vxho1jwKT
ULC5/eboEml8CoTaLTwMXqqCj4BsBoB8TWqs7IsiLD/hMtspG76nqI1PxL3rnlbsOGTQ2f6UISJE
SjL9lF2Jkjg2+ECk4M6xO9JcpGqSyjs8Fhe44xOMk5aM0TJSxqfWHm5X9T2iG1PTTLSXLnhDrMZH
7aKr7noRGp8mEdBj6TPUZshnfQlDrwg4ByMtpfLApfKvjepiZKDsaehgWVKmJU90+jH0Kt75wONC
lC8rLLLzy5/TOoEjWecqIVqw6U6U90t0DcDahB+Zb8UX20lnMsxaxGrgs2jZ8ZZ6CXuRHOH9WtyD
iNOM0kDn0Ffce6X4RcsHBytS65Ch7YE/2sR3owYUjHGzeihBwjK1wFLFMGHBiG81Agp6kTMvitSA
GuANf0cSdx0xO/8U38dqNuC68FUSNtp8JR7G+ynsZMUaJVQhYl6RX5h0jcbHU0pfY53dadJlxnLu
kVtJkk8CFQG7h5u9VtHglxJLyd9en225ZDLk13ZrQKYCUFNyCL5ff4UJ9r2bThjWcUZd7iIR7R3K
P2+nZgpjgXBqoxK6Ohu5R+P72/NcIVgmcdkHrS8nbrw5PUK7qCMJYDsVS/Czt/ycscNY6oBSHIBC
qlTfox6Sihgmyt03LfF5oePsm0h14M1vKOBU9pJd34q8sA3rE/F2/IpMcNear4gtRzSWnl/nRInZ
y4sG3t+XdGQwdrJXTpXkHlhLO27SkTWT7t2dGSOKY2LNsVupAdTlho7Pne49NsXCNGI70gX/Fo5b
eNxIp2FD4WFIxNo0j5t1HKeMqXvXml2soOnYdlyuf4w+IwT+v/Ee9QLFbcsegP1L17Qaf8bnAFdx
gMcL/EzqiL/ASmDBUciLWqjXOQBuiwe5DJ0jLqnd+Q1DiOKOkKcB7TPsWBJxTjvvvapURaa7ert2
OeaRwZYk8Sh5rU/XoiqWv2bD5k/MTPIK/3mdG8Yu1QrKI064WaZH6bBiVJJONEsuNfOhNQl3GOV6
ybO5LIWoHESzbqx4Dr0SrI+V12pcbnXnDCHEtX/f6Hz/edLmN9OqgrFh2SS7LM2kTLb7prRYVcXC
N/udSlTeG4XWl8qXUEwtdRvC+JuHDlq7yFMZGFBC70xlvY8myNV5VlIU4+ncsLkpL9d58tTp/8EK
d6/e9kG9+eWDsrwcmd+IAhGa49sypA0A8aiGE2BJt9VP8/E69aHmiXf0x2EGDsK1UOpYyylJ8HbV
1O6FOVGyyZvbTpEc3ogTfKRs64ST+oDi+PnIhcHt73aYu/q/IzTajgxNN+1JE3qF3b0gA8gyKpzh
vfNH4uDwE4XiQ8KfDuwgTaSsbvGUm1D+AgXE7FZg7ka0mwI2L3u2ggbCqnNxFA89lAsDKEV6e9FG
yj3tr8wlkdoVrhlMiPBgvxJJyLaCBxj8dqAyW8W8bILPZE0AsSo8MeKxLw6WKL5FsdfKsstwS/y+
IE14o/H3M3ON8cqMGIcJ17vdGjmT+wbU/N99WUQ1dTqGFwJJ8fj95LXKk84kdMI8KVuCykQnzgAu
3DQdBWBAfr8+k+4VqCW//gXkJ5JwYt3p1M3t92T1cqriCKlF6/7n7ZWHM60899SJxUHD09NfRyUp
kOAuR7MExHLoM+jZvf95eJGIenEFBQik0S6t5tvOLFYht3TnVQNh2u59J066cQE7Db2OuqN6rY95
DFfPjSaVpeORQvxjyH9eON9aKl+Rf/XuiT+SJA98sbnHtrHZrh7oCYGpmkEYJ5lx3TPrLR6qLjLf
PeYlSPtZWsPeaWOlFlo8SVSm+OMgdUFo4NHjYjMpODTw0xqUmDTNzwtEFTOdmkNmfcUU/V17TGTY
ihkvzT4P4sqLd00lPnMu4MZpxH1CN5GyDPu8tTRo0AkyEWhDnmDvQumKsIrDepA5iyhS+U1DsZ3F
VIdpcUlYCahQPInR2bOpkXpWv9wUXnhbMESvRjvHgJkmlz1ktYCtbgGKqdA0tcug4gHy67QK5oEM
lVamBN8FmOU+xVTO24j6NW9RITv4rPFtucSQHY7ShKwMhwmw4oGg85qocOw2R1VEvYMx13wsff6f
U47FSylWJVDbTw7sclu2QwGMn/xlIHmg4IhJFon09fFyvWvk/VqzXKJIUTMbeZAkQCKuMrMNPyS+
yyS0tkXKxRVFNWDmsUFcYjto96vWI9gE8pIkpxsUb+vvp0CRmOIw5IKtrisogteNe/boXrbrUz6Q
rwOVD0RN3qkzYt62T6Y25j6gJV/tkCCLFUZzN7CfYKLZ8FNc9K3afQkVkaOVNvL28MOec92oszH8
LWHFyB41DA4Ho541SFdiwuYk1NNu8nhmZSaudAcXLQcjD3V+IdT+dbJuteIERorGw5c3CZU39veW
aZhw5z1+J2oCBUrTTAekeDgq3WZzwW+sHW9PIT4v510Rd17nB45DXkUxaEh31SfVCwQ4/sfClx8v
WGZy4iu4Rv5Yp5/Ik5BDs8YMicCCrCVNxIMOyf4rjYvZdoS/Naw3uT1fJLVlNOi9UgqdPPFmnJyi
U01XbFQBdBoNNOs3YplCYxhsUSxNQgZMDDizKtb7aB8vT5ZypNBR3JDWJ+7zhKrj/SpSqV8knEVl
P4BjKcVObvOHYB6nSHahX0MTfaK8VU8dxn01fjGqQWoamfpPdC75s6ewauA9S8rwOp3pEIIDYpOP
d4n+wPkz3ctAd51Bf3JI8w0CcrPsiBg6wRcmQ9pRqfhXwNKsUZ+8Czl5zK+0LNsQk+rL4sclE1Uz
hRKTVg0PZcf0JJlAPstBHWlJrzTaFFAi4ppJRX2H535/XIN+bJpCSnnzHMxAaC5d4W40R+aAbB98
+6A9G/vox3AUCOJFhcGZRI86jTKCv+rEbWWLXeySe2S24FNDWkIahqnm1UWohJF2XcBr+KwNHUMs
GxdNsBpZXoiTZPhAYFVewlYafxfV9FmsItNqy6cYcjLmGO1nb07bRJN1CcR8W7N3BeeKR3E8nOtY
cEV/Bkh0CMjGvxU+K9Kl+SePeqB11iaVx7sdRGyrfl64WUy95/rtw7qLSBPlD7iZZcf56Gmf300y
GnOFKnquQc9usO5WHnmLX5lYPHlsJWWS2eEfP24WYCoQt/zZZdOyI9pmN3AnZk58KjaoDN6zaeZe
mXplAKKIjN+auzqagTDwUoZqf6B5SQ6ikV7cnRnMm0TyoCPeWZx51NIe/0qFpLh4LQc1j51rDApi
FZ9ILD72p6HYSusJDXWjmdhv91v+Z/fxd3p6KCIuvqPbNZ+JojWALjcoNmoYiwp8cBUftQIZ0AjG
zWB9g/j7L8KmuMwj3UCDAzBjKiud/W1yd3g+W34AKTs9YlZPL1ULhrlvogY7rBAX4zZa8H1Kjag4
ogkTX5RlOX9BCttubhggimtHZZWpw0Fsv5kuHVdLdIjTnSFB5DfjyErrdvr+OsgPmhKmuEY4udW5
qVeG3Ytbj1VlwGJE148zIB9CS/2pPR8ECdoKZXOc0C3ZL06R/oqY8eSIR385M4whytRBYh60g/PZ
CCMNXlpRBhXloI4tt83M4aBWfs8fYpDYQ+AQs3xpvT4DWXtzakc0fSH42zwk28ZX7KovVqvJsguV
ZmYfsffKi0WB4JUGj+KLYohNUzt+ItKzPZxLfBWVakMV4rzmjuu8DwLvjEsMKLH7v+qeK+OaCnSs
aQP7t98nzjBgrmTKZQPa4qPxcVXBKu3sMgUnleQlQysdOCIPKrtT2wNl8g3GEma6J8QyKlIdcVA/
wLbk9mC3Qk6aVBYlp6qzCghrcrzE+BRdVmOQcy/+9LPqYjWN5soDt0ulWIWjpPlFbQPlmaWEGrQ3
nezWJNgw5zySn93pRF2zNTf6CcbWJtoOhkhxckITNKJKbpRETR9ntvtTRnyuV4O2fNYe8eIF+dBE
NuJYfZm/baSVSBF2mOXxmpveN8mrCERKbaJz4Y3VyYDwSH9tYFAglTyYdv6apBAMzROnHJ362+sb
aXoV+sRNP+fpyLoCISMDdexLNxO+wDhJ9BejHu9hTJKxFt1PuvJzfKakReH1stQe69kN3NEowCjr
aYF25XCpisbd038bHe7Ftr0/AnVbkGpleJ+g6lfBfWVxxy1PFPafJwqPd/1zEemU63VmuM0HEVNl
JQ+hE4XZctEpwSenQEE20EpPacG8+kXHYjlNqOTAkvg5opl6l0NgsRITKgRCav7i29dAwhRjZ/fe
eiwrfPywo6eJ2bVGo62B3ixgYf/Oq6w5InGFphP7ZNy3lxIjWzXVaoeORHxOmslTF2NhyRNVxBko
nFEuRP6wP5VAUCUn8WNMeBK5kzhCq+DR3ZQVC1K3kYCONwqQa4qC5bPbJLdKKj5LCkzgErCbu8Uc
6Ja86b/3cNS702jZt36eQVGTE3XcAsfyqvq+aD8Y2Vyz/8Or6hvip97Vg30/NM0jLgMXYOM+Du7X
YxU3qnhnm13GKuaq+EOYmhs0R5DqDUZDXr3tizFTMQ5Ee7NzZJRN7gUSktBWcJBYik9GbvKlESNl
I8bXsi6DhwmtxtXp/j5SLtZiLvtxEKFGXGTGizz521Df1o9X8dwDUsKodc0mmOpkdy+vg/Hv1tlp
OZPPa1oYhhjENDuC0xm0JB3r2okoU3Xcgm8gXIEjBloBnGc1eYb/Ua4/v6qTClArXiBNWqYgpnib
rlpe0FR/us9PuqXCCv7LO49DzS/ZZ61/hhBXqqWA4tXiCe6CTxojkyOJZxGDSwJUC1HUQTtTM0+/
9fnRkEbvYHVsiq1NEyuC+ECq9IEl0K9Q6h2YMMvLWPAgS2eKlx80hpXq0Qk7uhtF9ZB/AvcTYfsJ
XB/QZ7rIA6/xq0RVFBLwfYmReoSVukWJzQhrn92RaoDJNWFl0v02Oyj4wQFjemJd/0wJsDV962EI
XCq2vPc8v1k3jiz4CIPTPg477/SAfO8w3c8Cdlk01w+XCvNYoJesdoQv/H7cFPwp08asYm/LV8xW
/MK/xU21BsFGULS3yPqQUwSqWqf6ZRGaOWbCWjfhdPSK/hopfeKhov2ABC3Rx+k5IQfeoOTWLZkG
jPVbLmwpU93pb3OSCg/WF3Ymv4/KmqoEp0OIj4o29EHg8htndFGCwgmqtqfGwBzBttmwCFO8xHad
Lq2O1lK79aiD0B0E3e3SRACCwQZD+g+fwCZHNeBxn6/3Ez0ZGNZlWsIhjJ4wKrrUQSaFPjhWdxVQ
gqhRC0SJ4fpPcnABJQqa20JYq15coxwWp8QHFrQnzDcWVL7T8egLJ6d07Zo8Zlfls/o29YvFNHDn
tz4mRLLYRN5cTyPpv5be5a47OGvUPVxaH2tI17iNsHRBnUQMcVVtGCSWmK6pJ64+aACAshYHaT2P
Wmvnw8AWN7nSXG30jyi2mQ62+VPv846w9EciTnlOrOg8vhkDuswEjBTMI4pOcxKlKgjPNMP9p6jo
yzsZVV1n4pLeWWntwEPCnQcdxGqC/YBc5/Mx98pAj4mbPLDAcy1uRcGbDI6NJNB6DgzqKq3I1jwm
heaQysAoH2P1AcToWAIdOFZwNSFGN9RVYaOUqn5x1/RUwUxUI4j1A45WjWV0RZCXa7kvqIzRtNF7
Ph7RjUsWzsNNEtodg9rm7kiqjm7G3fnmolcR7xQ/0L0Jo78nlxCVWuO7XuN7TN5XgHZLKQuwk3TX
cIa1MysJTQ+fHf7U2megHE1uGw7JgTPtInJ8vHRlO4n7OevVrfvgppfS0Il3Ts/xA8RZGINji0Zl
ZAkyeqH6uml51dMpyVmm8NBLmu7pPy+FmTin7oE24wEurwYtPTHTyjeMaqFKKzvXeK4RvODQ9iYp
ONibroY+afcDV0XJyT+l8aHzfasEqwEoyNSwkEbhmhDPKhtKuQr/Y3D3vsNBYLBzFCPiUW4IeIRV
reN4+5+8UutunNKkzOaLqhuCJZwAroMc8yyRSbctt/wMI8D8SvNksfTj+w1ROwraQSgdScRXsM77
oyMtoA54Q40U0l/6ZIKQeAdWobIzy/FYbyr7j+lMjlqX3o6cIffM5kZ9puTvlnwXLC6g9sj1Pno2
axvVkWWdBtzIITihwlrCuFMB6fFU5L8NLCxedfOMVaj4/D/urWGl4e15seeZNgzb03nJc4I+PUll
9x0TK00NYQLMAKhOXEDWS0JnVjaGginZHeFC8VyLPYwOi1d14oDi1Fuo03NlvEReVc0OS2BJMJPU
FjKWGWD51+683naJnrODwkDpXQ1QNbpyZsbtxYHvgBCcaktacbCiUWuiFDKgaHFrVqotXrENG2FU
9bMxIDn/S+HGS9pzoepRlBq64fLdk7qz7g1zz63i2C2oSvWeSiA25/HFb8M1IGSybpntZ3r/fIgV
Y8GOVbbBk8X/CwcVR1Fg5Sy9XvpqEcuhgcf4ZtxR/2iRv5HrZ8mNO24jgKHL3e9HWajA1Ynq73IP
UcYJJlZoICoge8oklu3INcG2e297KLnXAuopYdGCk1wN0I17CA0lRdRFxosDY146kTYRUjoJ6s6d
xveMRfrGEIB0laGnBCCzM7P81Btixcg8bnYFLSLBzyRXKs6UEahl2fubHeNF/9gBjeW4oxq+2qsc
cOkQFu6DUeo+RNkcMYb5SInyV7QM7WBvJePgbYeZ7MY/jIZzwUXfxm8rocSbN0A3XaCR9YhbbeH9
1eobqFo5BlQGlARrdxJNPTzWU/m7JCKkprgyqcTSLif4bvMjopbR+ZS4ouKtPKIb8hWWVusJ5h1q
D/7I9vEBohFQlRGGQGuMuKYZ/rMtv4HxWaLjh3+2vWgG4GOqT8wvWAZxwvXOjNjBXWwbia25IJbY
CdycZhZozKaMcTBYsGM2I/CFiNL754QrEmumWwsAwTJCb0cwiH9Uhfq1dXh6EUk3IvZZd3Qgp6VX
hcQQVP1XC/cqX5nlKOvEiJtoienzSMVT9uuk1SXNycB0od3ZJbJGbaXYHSyG5aA4xP9TXDEs7nbA
CBSp6XqUKxmSRUvLZTzd++KHrHWxA17pxw2zEH98zEfkiY6vW2Fo/9DqObi+a6hPn0LNdnrC4dAp
42Bxp15HJOqq0LBtyRJ6+m+IXO/jpu+3Bk89poXajgKmOeAMzMc2KNRqwwgVHle4XnEjtY6kgvNb
pGhXX9hKnsBP5ksD17e9/zFcLdtUBe+DsvLcn9+xZ58nxOEBvRLZj16pjMqKjxOFFPjh1VNhMXrI
GJkxDDwdA8N1m6zZwlDGpun5nnuVsoXG4bveBqZIOGIIp9b1JNqREuwV6QKjK2uKAAmDr66XiWIP
PWZuOc3XNMAlBCuvv/FKTo7Ag1Frk/F93mekyl1vsLPE8QlyWLi6NTrvJITXWuY6ijEzXEdO0QoC
Dz4vqPe9uHVMTB0N+J+FK3wR+Ly4q3xt4GSISK7eXZYFWYvRqJ9yGV8fFfcQ535bFsWnPVgzdFWv
oENMXn3EvxwxwzgQK2WlptzLVxHZZIOB981gNrh69NMAlt8eblLvFpJqKxv6A52IriZOemIdp/0J
Xv3LTX1lyjp9Q9r9tGS1MRKvPgqCEIRFjjoTf/7NVcqXfJqAt19uKBT4SeLHpSFb4WHyrIbMxgay
0DE2JAMBticy1VrXE+YkyDUw3q6nQBpBihlmm6rKcKyka7eoLoGB3wuP9ypGkGPDHxBWnjJa/26/
OxFQeoROg4zAJaw6M5Nlm5b5t6K/Mu3k0YGnjRLU7T6OEckJIqwLQmRnjz0DBPW7LU2HyRbkYEW+
HsTJryjcdJu1/fuYPe1V2/1duRU+XojUOBQKjK+QLqTcTjaW9W+nvTeP2FAFpCCrlAtOQatmhloX
2t8uI3MoUL1RWvieWSNH8W/msVYP7OHdh0w19LcykPOFxAovoxFWH6aQva0PYjtBCAShLu7zzEPM
QfULcIcYFxv9Jrd/cy8WFWp+X5cli6oGlWnX6Rzt6fd5Eo3GdYxnAOY7xZIFyjpaXUSLDk+GA09p
HFMuvuXO+temEdmiOCpe5Jf5Eym5tfjD9ND/IIratTKK5Tg9CWOmzma4xE8SwEkchOnD0tfEM73g
eVPuQ1g1xTKjYKRMtvshVG5rwXh17YbxKPT9S42QRo2YjDFajk0JXK+INA6ZFIWxSYngJ1O5qTxa
iKBLUfY/GMTsjslbmBm6rNRadNMSEAwPJf4gPKP2qoU1s4wa75Prl+QDd4c7FtX1oMiSPttH9Q//
21X5/ETqmyn6h9+iEpL9R94U004EpGQiCI+sWGSFKJiJQi7R12EUCDbWftjw+yYe5xeZOjDi1Yjn
nlZGG4In0fbUwNTi9LeoCw3t89D0qAzHD7h+HlBlvOTqUqoyB4wmtx2MH4yPMmLBNhgVtoe8TOf3
vZsVbDu6PLnmgdL3HCDclfINHjAD9Po4SoKPkHAStK7UCM3Fw4N0XJ4DzYKJ4ur64oDZ4AlmNGzE
OpG9Nffl5JadXwFk8bWodx6UGrM0Qxumc7alMtG+iEC0KcvGm5NeC4uKDFUEhUycywyHKVikFzFs
yPDDOgftoWYYAlgxW5b6v1GOQRrpGDJ63KTwQPITmvTZGeR5zp+up75i9tlZ41/5D44BGYobcBLU
keRWq8Ie8hyTNSHCMbTXiv3IaTeebtdS9pJOo7CH95+yvQg2gTzyguO0e5E6N8mFhTBKo7sR7p7Z
S78QbSohP964P21DjtlwBqc8udsW2YekgXEPgD2RymbOU9ismtV80sddllgqwuZb4pw6yE7XgUcY
dy2c6kPVPyg27YduKWcdls+VLZHoVUtS3vzHdszqW7VvH6h+hVz231JUU8sOqh3dx2Rs+naUlkOE
YArOoLjLNRIHSia8JbcKEXKFnqGglpu8uCHCw1T7NK9n/yOftwwBBwhWEeDHccGr+hucorpV7coS
Sw3ZPH5yVrVxtsFpJ36vwNo0qOXtWPMb6fu3dGNlEEFx7Bjb+ZVuBo8ChCtlfuOcjhErBfVFhekL
qEMnCxdUVNvF8VDNWj3GM+qu9i4csis1NCvCkswpYVmat1h0rYec4KuHTV+cQ8dAedGGqexJbJ8F
Eedp7RnFXIdgrBFjOPDX7gsFoas/2NkrItoobggXdB4gPkOKippMa5+ylKUaWBEvPZ9U6v4HdGXn
gVP8o3qvlzOjfBedsxJ5JkBJ8qembYka+9BxlorPzkXm+GeNHAq7mYusi7e9wFKej5zS8RzgtTjX
QMnpqMPlckqvyymKOoPdOSpYmK5wTL5sfyfgxI6fEqQ3+Ws46vktS1YjOB0DJTHFPXUPqh91iOaG
i11e1Ce7+f1tIGABCSicFxW5cmagSDjBN9IdkLtyL5xoro/bWjn8LpLS3Gv3YVW+rNbJ5rNgAO9/
CG1fEgtK3FJnpsz9CblFy6/ZpJ0yoZ5MisaLwdnHTXS5Al20/uFcs3OYjOZgy7ql+p+huDt754vk
5c/wStQ5vUsl+UWrqlcKb5lMnoPtejXtv4t6DQIwGu4L5IA4OBYsCMxbmT5kDRM92WSTP/dmb+f+
WK2BtgzZclnYbMzxoi0aLL62LK3UcYOK4HyngGC0EMXfbMUKT/ogL4B+nXlllCeT1OabI9Ydyi2l
VhL1TihDHpBuKANtSTsQnOKfvcnnzTt78O1XgB6IokUOljPLBEZZKJ2ORCr9nnUO5XVM/VsRjnH5
IgdFNXwf8oVYhzfzNEkEHaWBLklo8tZ5bZsERNSeofLC3ZL4rO806eI3wjyBGrahqFNQ/5qCF4aR
KeBtpVCw/iofBy0vV4gibOwqrC34+oxnpXjmCuDCB9xdoIy6zpjEDVNS3WAmAol9wvr26WLqQZAC
QYKpas1k5qIEAETjTJjq3ERpmBG6OaKH5FiHRKi8Zc8m4n1XvLZ1PpWl7xQRIrL4D5Nfz7C40hmX
A7m5ITpeVgxZf5xMjkuedz0c2hOkA8hQWJ8BIugWyia/KZldp7OsNiurFIcuTTdfgYI5fhrWyRKE
qNxp2idf8SGjbUR31OJmCfazBbfDbq/RZjOo2W6WjNZvmQeDsZFbuXB1/yadhXgHa5iScebwgqWY
LijabwJzb9axMcmD7EU/L0XDSEF7taCoGjl+Ri3W6k4cC3ztb/AdgAFwTVaqHfy6MQsleQZkZ+zq
WCc8M4AJbEYnljMIV9WtomvrUGGfZPLDiu6P5qxy0h0RTnpLZ8HHbTAOBU8lIKgMdwvaCir8t6FI
NV5BXWr8U09z5EjI+h2fKQha9JPP+lJwY7T9VuZmiBemmiQaZ6k6nG6YhXEPK+JG2fzr8EMIJh5l
plnCTTjDMekY6xuLV/Vx9LmRuDhr2IWQ7reLD6uGlUepx9s68oMjXD6zwXr585ICpYb3Z+yOwB9g
FeE77e9caRtYVN9N2v0QLYno3X9fcqkS3Qh8yreouc8xL8jAsTIxlbDIMNWSZToxKOStvdiD+/ZJ
5dXwY0R8zekCtJZBnVhaEUACUeMn76lKnd7U3jSazPKebIg4a8CreasLwmz/8gMi44gB4HYGmWNa
0y61iBhvQSMaoIkb8WYxQainfBAnvkhaGAXscpz5T5MnyjcYOmt53qVTOU15PWZZ5fe+SedFGnMd
rycNhBT3Od74n24f+SmtKuBH3fVzpxS62yhQVzZ9omTd8qAN7ugtbNY2dGxLoL9lwl/tGrkThkHv
CkxL578QPoOkLlNZL52ElzdT5TtkdFmW25xbV+a6zw8dVAv/Sh2lXpzea+GNaYYJ7DF+DdNuJMeX
/goEjxfHZF3eALCIZfyXLdFJrAIkWgPOvMfZGkSKddtPfD7qJC7HApmpQ+hSN/cDPDj3fs+dvgQM
H/q1FF+qud4ckex+28l8S12/xd4jJTdR8IFZw2atQmxztWVsWXdzs+cWx5UyO6LlhGOTOv5r9NTx
5/MeMoyt5Kavr2IHZBw/cH3GF2bI+6XmLiU0fJLUmpqGFGQRTknFUPsI0ZIPD1oe3knKUfE4zY6K
0kJnX2dxknPkDXefRu9uV288H6TYepT6aHk13+0g140Q40P6WA7I/Eb2LgDXFYz+N7J8MWsh8o9h
x+hOhyMbeWeSyQpDS7pXb8AYNhldJ0dlMxAhWhqdnTV+ftc2mep9f3kklDrl/RAEAQDINzeajfzI
mfmKoauutkqHyBrxiVAEqLS3y4auUmvmfO4Bs+CKnaZSu2gi9irhH9xm7A7rDYpjdmPOo5NY+ZEC
e+PUMG5gIXgzpnmYbqqvo3z8mUfB7pVTl3o238s9QSBg7uaTSiIizliEGQNyLlOS7PwzEJR8VDlX
tiw74bm/yNM2M2wqvGaxZNZNmp4QTZgI7PCuGg/F3vTxgQzG8FD0eZ2aGJggMZHbzW6C+DpN06cC
lk++2S4fR9RWqDntMWYiLPhLV1MaOQ11F0F7rtvb6qfjcPZIdy1jrHJT52tV1F4mY6M7m11WHm1r
4EnKCMzreJFt+DvB5+Hu02S1PZ0aNni1snM6HF/A/S2JW/YHQBt6wJY/4ezFA9y/GkXjloSjd4Nw
iON6Epf4zp9iFT/URmKVdpJWTAfBUOV5Q4+YwN+ZeQ7Ud5NqC6VbzU+3pRI0NSNDqoGz6m4hoQBu
194qht9K0t04aA3cciLqYaLwsn3W1soU8ShZY9NvhvNp0a8Eqv1AgbmNLuFQvWUd7uZE8yk3t1FW
RfNzAxY5AKS0xwatt9RbuVDnBmoQeuD5xKoBQHLbHd4CQH/ps9c1o6vKFd+1UwAGo+jxCwr4Oosb
vx2MYyWhAF63ndaKWv6rlL4DNfL1WCWN/vbDXnZivr394mOapEV7VXr/7kXHGQiSLinSfc6kT0H5
xuXwLOydMvP1WJqhZmeayRP61J46eqIMqsrF/9GVMkTBe5pib5f3SQ+VYXY3Brru7X59dWmzGXQd
86JdqvQxFkk0lu1y4+4pSKG4H2BNPVmEGC4rt9KdSRCLUCUDFJKeVuN1MUy5IH/BacADRRGq/MSR
jYoSgG+FggwUDXBSove3WCJNYT983VMaQACBt6fUgYn6l1E0YeSwN/RE3prYN/cungz83sPdyqyY
H87NGWS5P3jZtesA3XlNLhe0w1VXlqkElOKYjjuWc0faFrsUljFZfJxgBiZIQdBzSOaPUJPX2oGs
yaH6qi0C6Nenajd0bPallpcxrVrMFvuuze5aYmY+BPAiAX+sXQzmepUzjNf2swVizi/fMlTzfB5L
kTwWJy0nqaxZXr/ix9hv4tPHxZJVLcoATMz0KA1HT4eAmypNCuqDphOQ8NCsjjIwb8TGgf85uTrq
RJpufjK5R9PiaueCeMiEQAzH2t8RB+Bc1sxiUHAMT0ww+ALCc5/iG8zxfV9RqSnGFrrdrDbTKlX4
sAT7KQuYbFQPPnK+TrxW21VJWNb3uRjl1X3ePmBlxvO+tmaxbBkDSzLhYLSaN4Ye2hgy2CLYX70y
J2RxfelDQRtWGzo9BztyLEd7EGRxVWQs8SoUjMUVJUnPiwIBJ6vi/MEg0817P7WloKfz9BAZVa/V
AWpu92z83RDdrliBN7NWc1vCcuWTFf71foJHbI4Q6R+l0Yuca2sD1B4wGvkJMBBhfLRICoWf2IzC
SQgPYyz3hXZGGNMXiujlK55cnc3Wl8OdEDWefSsfzFhQvC1jYjtcaT+QGdDfNyFBjfT7/fjrJIwZ
RThCzebUPFktfmodl9oLXjMCgYTcDJdDIPGzECMAPIRuZJLQo77iy+QlQVFnsHbu/i7+a+Jc3AHh
spkzeKlxaRUJBEbdUJUpYD3hOAXeJscXQ/qZhs/nx79PRPU3kFKOCe6TVZ9q0w73XTPsLP/EYZln
/xPkClD6xe7GJTjTauRSJSYBvmVqEvz7yh69DbUU+Soji+heD1w3DaEtZMPuJniUgjbR2RvbY2pV
579a0j9YXCZfa7g60nCtsHeH6gY9Sg8AZ2kDRcfVAxMIvgR7EhmyPc2Yvxj06UK8MlqK3VPPAGn1
9iey92Q7z4ZYzovZNJFnt/BuK0qJol3oI7TcrNuBDVHpe59oT5Y5jAoOyXe9H7iwzY0EquRgWC0e
1zdMvDZtkAOKfAGFCdzPfzlO5WcMBsyVm78cPZX82MgNgg7bx4v4Y2zExM8Pf3ZkIaiZRFlVL7lO
MiUMXm/ZLm3oRWbcQmpYGZ68i8dVWS50/Xvq69cw0X7fcpjDdzPup5z9NUfUjWi4ogtkxndoecXz
6h4MXRpY2BzcG7Vhinow3oHymWmw5fHRlEsIr0ONO+Nycc398ZTQoLl6vFJ3uE5GwfAS6kHS89mM
OJzSmCQeEVf8phxesRe3cbmaCk9JkF/+Ev5rfNCPwseUwKlWUlX/2qQ4jQ0o8XVWJ/WReh47Uv1/
Q4mWOZyoE5pt6zuzi2B4NEJmkdU84q6L9t2GLMkvf5xndbGu0sa9eXFUTJwKya5cy0sYW0bvfThq
is/PCZrKLGJJEZyGUeOE6mV8PM5NY/oRjiUi2jO00s/iXXvkfxcn+L4x31ZmA+2rNelj6Suu8FG/
lln4ptET2F0KcsK0Rb2TNFnrGlZchtQW9CrfGWp9V/am+3j6RW2F/G4cSCwL/dmvJmcEh8AIGM5x
r/Br70FuZt54v7VhQwNaRl+iWfuC3v8TcJzU+Kzr2iQFJNLKdK+42XfZR8h9JTmxs3prMLcKYQMv
zDJhdv5PmAYSJresTo5Ue8ReHz9ul4R7tZYYN4BUmvL2mmIKttmQAfza7WE0eYX03B8odWzWrgQZ
rYCKBuL4p7p8Dik1N/+R6agjyBn3/68rZVEbS4MRlsVFx77iRvKlEt9gAq1kbFMPkMqyaltBizOX
GFLW/3pQdLt5S+/Z2OX/oGdl9JyfFs6XDFPESNaQ0IcFSn70m/xYRtRe6Y+y2CGUPBQw1jSN/NhR
Yd2O3DFXOqrrUOzF8ksq0TqbqWfusL1KudpxMd+qzqS1eHlVkLhcJfsLetk7lPnJlCfR0oysVta8
36STrYnl4g/Pjl1g2t7PXt8SXf1i2GGgNWlHGnNQTWKB1afxTF6WxZbhmRtr6/WRRGgeMkaOE78n
BNKsQLVpB0kSxlfCNDeZNMOSdnmQu2XkMUAF2FaovZbDRMx7VhAyXHsy+4ekKQOdIjFdhaC6CY+1
52i8PUJykd8EnRzOWVJZfBJ9DMWPwwFDUzyUxPx8hYOxpyHfpk+6jkt93xw7kzPFg/QntZCLxs8+
gHznlP8kPN3xzvN1/Wo7QzI6Tf829qY0Sft+O8X38NhyovokkBCZ+RppFBdf3sD3NPJEsF/jA5v4
Mk4fn1kepg28VWehOusnuHaeCJRkDttBNbyzZLDlvA0Xsmrpw8vwbjojHgqLkme6zatRoFU/JEZu
n+s9TFdTucAYbTdO/kqkhmW5EG1oOtZH211bLQQmQu626u4yZ1juGECH2vSTe5j4wh2p52wLQWEd
7QHTVUFBWGbDpziaDK7B8DsNAo5LRrV5p4xDhwjVYzd2gqTIzD5ypM0x5o7v1xaxT9bXN+2Wo7ZW
cXm3mEeaR0fpQYZk5w9AsPV9yDqa3bhAPRs2fHmb5ef8gsdERPJhl1ic7zmqvpBm1mzS8GPUy8td
HdO73uMPPVXS0I88NlYeixxzj51AZm6eFzWRDDy6bm5QXMCt90aBZ2eIi+vZdiftjrSugLlkJmBC
Vcc1qBVQM9guklDirKBdqVSQSZkNG9xOFYmp3D3quLszGlp/QHpNInS2JqsTb599r/FnLGYKyu9p
vdU9570Z+/STA7T1cZLuo1IkZ3hVxz/4441BtNBdoe4u4Oz3pjfHEeS28Az8bljMRrKdwLNVW/ZX
3WvWcNaaoSAgRIix4+LJig50iOs9cg/9hpSAF0OVFayTNEsprMYaCJT9Vzw2ATW7msK0BE3X7FkN
jl4J5EJZ732ybmQdCXAiVZlAtvdejrIZX23bvGnqq0+X2iAw6ee1S4+aJD/1jpn74xwfo72pFJXc
h6VHDeHxASLITnVkfx3mRSOdkABKug2L/tf8XH0haNtwE4ts0FmUMBNk/RaoTGY42lNpcdC4v0Kc
RpCa0X41Pf93jTW8DxF5AhSNrBRkCBAA9ftaOz3qJGHLqYNzDnyNLRs2LDAvDCGU0iJAUSksDHrf
Kp0uRgfNRlgkFeJJpngYAQZb+mBAUoCDGhnQXWpUWPtH3N2gOdtSOruRBHEpSR9hO0Z9+Sp9b4Ow
v/cGuwo+F2cHUcQOruiKdWiuWBa0zADiZ4ed35nAmkhXw+rokxdr+RO1jrtMnmD/jE3Q5O3RGTIm
ZqELm/Ad58dgpNeM8+aou392QKLqRjzxD2PWpJlXrK8S0/j0lFGPVeUXdB8frY//xSkonDXwxI6d
hpUNBLLGEm2xf3OkMCMSKR/kZsMNmnY9N2KJ6G1wc79p/Z/6QsMjHiHCKFRgxiXjOdR+KY1s1wn1
Jtvri47/2Vwxzfgacm+RF83ZmpO5q4DY5SSL8iFGdsbRaIbqfE5Qq4bnnK0ldYVbJx1DSMdoqStG
a2mo5IbCTDDaVzwX+Jaq+srU7dNdPgbnoeMws1qMBnPJyLM1OZEy5wympOkvax+z+ZSSX9GrWWTK
3imx0N319mb+THNmkQbGl2ClC/WoCnebduOCHY3Ri0cCKymXyukJDKx3BAF/cCkAmV1H2l3HOgBM
XW0/1mmyBcXNuTq9szq3GuT6sBxrSpqjbhdMe7I3cC7w2XAJ4aRN7E2pikB5sLdICGgnhS1bFo+S
Jun5mF39PxWb/PYcPtxTODm8IMmLqATsf3nHlxKC4UbLbi22ZHm/rGAyYX82/TXURlqUT0XKVJyZ
Gp0ofnKF/XY6ysvuVHM3YkUytpa9/Pf5uiygPDg9w89EsTdl7gd0ODRtxXaW5slrdybRwhWQa0WO
aUe3Sl5N+rCJj80fJPOXiIDX0Rl6vmpvu/rtZsiLfc5YYzsVTGJ3usll730XJCSQmkLsPHT1dNJs
yu5mWm+QAlcRlxzauzJ4ibn8ah26wd9ridvNKfKTbcm5gkHPGO1EoXipZyPaalgI0BCdLT8MtENx
b5SrT5FbBYT7zs+T495mZAyEDmnCXHLr05iKDVdY/TSdoDQs0qTh5B8iOClcyygwJMbyspFl9WgZ
etZmnRKzR84OIIbsxIZzPjKv0VSZU1y73jons0zfZfhDwJv75m6QPQWK/SjWT+aalpNgrr6CxpwV
SeTLo0pAa6uDOdTnLv9QpKvZIYAE+zJVSAVj2iTium8YHmzVmDRZ9m+2QIbtPqL3VNtcaUVopdku
tdmsnZkStm+VwrEfdjzDorSYeD0m3231gQogjILVChZDWPrwvUFY+et2gLj9zSNGT6SLfpuhefps
uHoEd8GKkXNcdWEfsnGkPEuz5BwzjyEcCm18+oihxZX3uQq5ghZHiPoIqY/y3fext5bM5X1sx9+c
TQT+HnvIP+MwN4BVAHmqtxrYzIHMu9Y4gGz/trJvRMwHThYZ9b35NI7Bt704p0l7NFhInTLU+Vdw
B7JCjWmfM3wE+pnJ0enZDty/ao18nbCdpdW5R7zctxp3WXrsZ+PAKSaUxJHfiPIo6D/E5Va5W6Q3
I2uWcOTFlqXeFx589eNaR0Y0tCsPsspNhvIEBnk5goiNNarP7qnzqBLJfb0J1ki6uzR1Whq0CCFx
xkdzk/NGSti6DFVqHjMmPT1e49UvMpcWS9gNikJtR90VRGd4i93otR/mkApA2UQgsaDC79jtIlqU
JJ7NRYf40i2eVMFUd28bHgIrkvAZSImEG+tiLREp3qMzyt7LJKkHzTxX/hrthAhvYXBFtPoHNGKb
uYq6gBop/9fL9wdVyC+ne6ah5nU+9w2aZb3xcAUkOR36qA4Zy+4i7hJGchMs7zL6VNxGlmjmD9zC
ovHioQUab6QJsjaGOXHkDkFbNk9DhXYby8OxsluE0Kza/TACcsdlH/7KCiZ61vOM0zlQaAibSGvG
pHlzwC20xEDR/07hEmpTdGebaGxm1NmQXvCtdpUUf52y81fP6GZ5T4MrQNexZi+VVda4Te99ELO+
yUdKUUDJ5csNTVra5DRAycDH2wvcWGTeVaZys/xGxyXjKNl9AL66SHRiJUowwY1wqQwDMLU0AZov
OZ+nOMvTPVKx2+uuoE26z/xJzsNs3q2EJN3MpmLyDnBkgbQrmWRwSU07Z59h73cvTcasvYadEoti
pFPxZ/NdPg8zY7FBugrEjF4aDxcRBsp9xFrBB9urlaTTuQTADJYR1yxuy4U8dxj1Y7HTX0dRvBQM
tHn5gXK5jRY3ZRUuOcrWcQ60At6No+Ro0EB7KzKkVENQTwJ5i6OEtyZ1PqDd1K5+Zz3Z+L79pfLL
2vb8+84E8JViPaqva42urQO56H1IQeZisP3lWU5ZxLJqMudoBEoJ/ZF6WRSYtI2XDK/gm/pcC9Vd
lAYIdb5s8uBYpp+6MUOdyd6NJaGlEVVrkxnHJ5AuiuAf0xFkthrxvjQR8VlgJB84cnTJhdweqV5M
BfoX3AD2s5rDrQWvkGEtBshjgaPMXBIxk32DeLHIRdYeavk45GXglRUuPwEBipoftYUK90vkRYi1
oBpgdGCm/EgACVInOwXpqgSd5V3uHecMaxTE3zRgzuYddlhBKHxEMb4YKuQEl48v5HegaCX97LKO
J9X02RN1FWfCq8QRJi0qiwvAXVAyVs1edSm+/u7q0TihHK7QZ1HrAdw1wFMy45yxQj/XFDpJwO2n
f1J3XA+UZZJn9UAN55f0K+lSltAOxutK/w6NoZYeq7mm3VODn70eFxm87eZZ+lqanz7HTqtP2H1L
CCY5eLNGqwoPjJFXwMogDjuwO2tXiZWaEC0qasmZZ4Zq9sairx4smUYbd7gz2niMhEKdDlYmuIGb
meQTKpsEmpnL2DqikWQ7e25YCCfQGuCQHEmX2DF0zgYXyEpTAnE24ZyBRae4+Dy14ngyFYfZHK4e
EDE1jL/hp+gJmmU0fVLohxLjzr4A9Yk8TuNh/Wc1+OHqTFe0hB/3YSE2hrlxcGsdeVbuKw/NEvfs
SdvsYLShwVFKp+2W6Sc/kMocBPzILs3nxzLePE/Hw6C5AKailLZtjvyi7O1E4obZ34WIw5xPfD9+
eF7xnmLBXLyXKcrjTHt3sZe9vLCKMlLuLvs3GSHb1TmMmd5dORSTemGaena2i4A6ONIkpeK10hTt
1HXfe7N/Lg52zCIigiOVqjeh9klPMwe+zPJiZy7G8q63n3jCR0x6BTi1TIemVnvFBVg+j+8jkb3P
Gr7l4dgi+A1n61guwPIt6u4/gvQC5WovLORthR1YfbrrYLo1VHiBTNCqi8ZIFov0v9BpxmCzBnQr
K/CfNTpxe8HVBodtPCnCIg/KQdBTJqVDOWIXJBGPIZhVI5RvWh6GDDBQsrFpwIVbn52roNi2tnpL
WIHH97yM/xP1JGAAHQhTJTbd5vHdDjjC/9ckJUCt9G66ZvsFMEP/1aeV/1C8/Chnbg8NLttk7Wuy
rBpq5fLrKwmEa2LvI/7XsZnb658uDbjWdNEKgi8YDPbIfWxr86FftRsDRjVTsaIhRSoKwuGBXYCV
JSEfhocY4Nooe73cXUWBEX1FH6g6IdSacUbb72u4UR3V0Zvwa2HNUfRg8FHyX0XZFMYqjsCr9aW+
HRP4xCrRoOC0GWSeLJX2Tua61vb4BCVKxUKRG/FJ8R4whRrCu4yudT00d+nCXzcqynHo8L3GUd5j
77haf6EGrJ5O1DFhTsr6AHnNKKK4BkKGH3S951Bu9+nPI11zDH00zG/Qhu3USxCHgyBonzESmu+W
bLQ7qkrjwb585h2sK/PHLViFyuc+1Fe+oEpGS2xCBLJbmOOs8qdp1uveinvdqvQPRS8pVzIcbYwO
nR2mY4IpdR0TYPD8Wtv1VndPVdk+9G8UwfcpiHodwNR+ynCiDTKdYQkftkCYouko3M6rWY+mFbWf
rjBWBkQBoJFunivU1xbvwErvn7cTjHWM+bcbx/ENMXZNGC9NJGP2ZFwKVqvBrD5ZLAz9YjvJTk3+
Xi4+uEx9xcF5QeU1RjvIYRmWXeLxvyeufLMakMxJ2igMFHypM/7wSQEivETJVqWL2jxv6XtDK0mr
BAiZk+BocKA+3n8KyaCKVLpLNYPPiRNG00QSOjVS24uexxoArYsvgyJPWdhtHZ/pKpzBWJO0aeZI
1qTpr50GkwEzJPxFXve+V8SsnkE9I6Arjk/kQowBLtukSXfwXAD1VsJmjVM5ID2+mvT34Lor56EX
lrPAbqblsEXvokx3VDhYkfN7h1NukOMoav7JiUFtclnYMNgoMubcrMXmydMQCd3wKW/MLQiF8vl0
Jy+fpHDl4j5CKvszbqcx+TzVgbDD37nyTkMJrPIc72JV7ohilS2j/Y8Vg5f8iQYNamJ8+DPvk/xu
o1LL2aFOjGSRnVH/4L7a4OfCsJhxA2ErFuLepSnl6r7jwMhkd8isCrkaFHrGUFXXQZ9zqPXphbdZ
DZ742j7eP10Xu4ALsW7MQQOzb82j6F1kGsyag0aHgXQfGSFBpLv4i1N9ClepVjov1bkhBWOVmKKv
42K0bekBNV1xTOUdDDPqNSLrmKXDBNFcb5q3PlFE4VYvmPgaiBfQRRqLzbKmN+Naerp6aevDbDj1
urRsixp9SheEzwVReCwhXgnIKu05zzfdQXh2yWfpd0m0pmd/TRGshn77+COZWwGzEVDzdmNQPoSu
kM4ujMGeaa29GU6805D3pcom/T69y9ldjXrcbOjFVG1PWdcNXEEVliOO8Ky41jKR8gdF712qHlon
QDGwTOLkN+qzXJnlHPg5L3amQ5LPi8VtyrLrrCJLeOuCMhkuN8xxuJHmyM9cu8ecIE19F7/YNWTw
xPr2hG4r4tzIuhfmi6yqy6p+Qd2LnQHjqi0Vlz/iSr31RchOFG34w/e7vQ6MW+6joOiwWyiRDpNN
0oDZ2ekhDZaM91M9NLZ6MeFetIFR8Uk2Kbske8XhjA5TqLr0GwgHoibmRTNpZm40gl2Kx1tw7Kph
Yge05Q9wMZT46xvadyN0rm0mlyGw0SsBpfXeVSPPM4BLOZ0tOmVt0Lwyo0fqHEoOs2XPeUgA2H0A
sEtm0o1oaDeYKYHuYWJrfZy5mYFNms42tU8WxSw7LBK/lALkVjTGm+LBYTTRWgGUx1wBbYjmdLT3
kGnGhiAoiFKuSIgoVQ764Qa0DdH74e46eY8cf7VXO2uTzqtbmUW9zQLVO4RAyJ5XyrVUxzACNhNv
+K81p6MIWPB3X5iwBdHrL8T6peoZaMHv0gfQ7utlFo0jJiQF4sZGRscIWMs3joTkWzn9vviSK2Bl
v0VMPWmQnQURc6bmtFdT3o21tG65rS+zotxSbH7R5vpuk5zE025lfxorFkp4jL3xECCzHbP7NROa
zSmgXFs09ueaWW6O/VlqUCLqbv3j8h6QUWmijHKRjTeGp7Lyi1mQn/HPMsWG4nzX6NJQuW5T90t1
eT0MzfpDa9hJKGlrNKGLY6x/AlnINVAv2Z1q2URs/DGXl5mEP2qDavFZqQWuQPH4OE6P0TWY+n9g
ZJDXBPrkW7vr5KqAdgzN72JR1zOWT/rvnx/IISBfnFUjKUQmxNw45tW5LnoMFMzqJ5USc4ueLX1Y
8+1QShNhJlbrWuCG3Rep6S8dXf0v8GZbtLl0QihCyjy68BzoVKsutD9V44XFQ1+uPieuy9Z/ExCi
aKT7iEnNiiA0PpvAIEH8sJllbt3hL7Xz273LS73O5p8+9LXNb/e3zImJ+BPI25B6/Uyh/9sc7EkY
EWEHxRdr8zYn8bcEaBMw6iN5pnX6E66D0gneBVZWa2vY+/0OOjHQefcKXvr4Nnoevz+i0noVdCRp
mh9mPY6hn2lPF81wywkKicTQJyFHDa7QOR8K314PcmRyYMfQH29R5qP6KvuPFh8R6f9w77RIivyG
FyCFYQCZnnsoq0xAKSwuKYFi8wUHvQygSF9onnfFzBu6vUJHRxvK9DWBfnsgMasZdjHPxRAeWgIi
qkurBplxzR77VHMWJHb35sZbEjljeZFexEfHmCkWeVJO1/9jeJ5hqySaQkHPcn+36yJX1djK8Zu3
tYKRIYV6RX0tfuBVMjSSU6xsH6cClF8SX9NyVgn5+upxw5kTFlP6qOhJXxD1JCdEkUGERjEr8Vpy
azNwU2UbkehnMlerTrCZjT2Sy2WM27drKZQ5849xLW9XFrLksZT9p3x7AEoMQ/QBsGW56i0JdAbb
gBa3/oXq1elVoPOcsRrTX/VqSPIzukzpEvTt4afZPMXTGSuB+APLJsIxRFsh4XTcsB3go4OXr8ID
5dKKEaJbE42HMqmnf+2S7y4h1ZA9EnrQL6Az0/cJ5IkSLcDut51ZxslmlMtQsbnVJI+hsWqC9sID
ycSqccPWPT3RSDmSemzus1pTO+25meEtHCHinmAyy0OI8BoWP4U5ohX+scGjk4ayOCoCAj1+g3Gg
57H2/OGCVtNStSwLESepm6Wo3sNYGkQ59r5NIl89AjboXv4CA8fo+5SbiFgjQASxn5cPgx2FYJMv
qbj/IMHIN7JgEE/RYg2jc5LIv8vK8hcDRvdQZkVdOuj4iamzFX1FCeIpMgjr9BzSmYicRn7CPt28
XO/bSieUP+btH69tUcxscU/VkEnuDVsKdjKndFaNYk5RS4IfIXfeO2ggCaL2pf5pywvSsbRmmsO6
GEC2Hc0yA8H1MsfxFaqR6qTFX1w3QmBqOjGHIoqgpuktSa38ETKH9YzK4zq2BRzRRcDtjD086N0t
+aOMuSN5wJqe8pCf/HXt0GQ2N6exMNHWRKoolfB6hgSwuXXQzT0dWePMk9qpm5atLyZPI3hbjUPC
M2g4Ut4RluTYLWsCWX3A7tBursavbeGZS/5G8lm7YBnQzhv9/7EPa7MxRlG9DAjNWtUzSr8u2juY
Xjaqp/6aQAmjDOJYbKweb1hKzuNt0tdiBFQIBzTFsblAudqOY1PWZGK5QKVD6KEMK0vEJqtiVWpO
AnG1Ho7tVLwsmIr/f9Rlo50D1lFhnRpHN9t2Kn8tIQLAZKIMJ565ZZklBxtO4QaqdctRe9zRYCjD
kPKG0H0F7usKoJz2dklHPo7y1h8HlHzL37G/elLW7cdTkKZkVkVhUbBrFysSBf7COwU0l/w0eTFc
uJDkp7QR81cwgp8F7xPxkg4HyPWYgCNVFtSEIa/vlCMaTBBsdnTi+K+tQKaaD6OUSBTJK1UkS8Gy
/YTroutRqS7SrCZXqP2GD/J39lZM5eqXie1swMnbJ8RFEW241XFhTzsdVl1j/M2vHikKiwmrWp4U
KztC4ox19I0cLvvZi4LadAFmMkPEiEp02PhCjmMMRaxwl8b+vK1hor/Nmz5wLTB+W+Bhui5duv71
AAd2I9Jf2fu5bxHQ6qoBWO7WEDPmgLXDg49PJR19b6LE8vA7aftWVCi7Sl6e4E/xwvKiMKRz7MtJ
d96eYWHGBLDOu9CbB8lQTOTq8cZnM3LiBWFs9htIzPuZ3UcqPRyFKMPSoWPhZ/ha9oCc6VrWNr8J
eD/iEnwLyH3IFOZ9kHm2cKL+d+TUt+CmIZJQvbUTvuBVvTq9MmFOHKbMrP5dVI+4Oh76xw1bk0VL
ohMyC3bTS9/b9bFP6/OFSrHGMORGKqPC/dYYxj0UvbfGqRSFQy82wAtJZEXcLSEMuRPWE3JoeUX/
kE7LBGpo+yxFf+3qFtpaynJm70A7fTcIaoEBx6R8I15dRedDiVVEeVp22C1a+Ijefvpzyv1qwTOD
rirBfBOxPScx8+llt8m8ZSaSTmMGAu1zkqrx466uKiAmscFWWP9SuoQL1axjBX+kl8GVQ06RBTi8
DqEkCSYS8inQBeXiCB1MrEphvlo+74tAaq48pPjTvPJkUILdEMVagSuiGxvaidGG2i0EXaVqYwwy
oVcM0vTGdR6c5y1zBjN5I3vnVaDjwc030zbI0CegchTgyU36OeYaNl4NCx+Vzc1oAID4cZL4GIRt
2Jh8hOBO0r9qyv4LwhKsWv8ygb2gjIT+hUzDucVVr5MVmvkOJ7PcW2DERhyA6E+J887dIfSPf6Gc
4tbFaDM4WeHgRyW4NLYvDuS1QCdi0cmqzNcYkI/mBahoWAmT2aLANkabwYrRCuqKuabHZXWGkrTn
rI1oU+mYaDjPACgF+lnGkSSYKD3d1cvkYsti6f6pmRTA9flJoJSogUzXDly8OGh+N+aQIq43QGlh
USCKGawuWUfu1ff8oeX2utyQDLx9csr7fCZInLVdmLRFsPUucPG7SBrqqYg3g+8os4sGL6Y+R1T7
f8Xg8/xdKqbvXdGSfXLUWWkRvWcdb8P7j95M7P+ZhbvZEb/mTAnEXMJo3ddT6RlJYuVZ10Kib27p
OXCv/W5LzVZ5phw9S6e0kWZrp8zxgTNIWlDH8Sukn814rElHxRk+pQwnKfHNEfYWY9qpQfa/l/EB
AHmffZ4bu1218O+TnOYYeFNz5od+bVIKAZMY3xoJh2Zz4YdrRgHstFRsihb/T8eJxI4N8bmIqhKo
O43aDx0D+8m2q1A76ATeFUuVLFbaQjJuxzqhy57HCqyDH6jsdlqmAPEle6BCg6dQK/+uaYchJwaC
G+Yjbd9HoK91orOyD2cn55dMgGEix40cxcxezGs14hd4bwXG5vNdqU5EExJa9UaDhDaxNjbGYIO/
giFDgEi20OEpSQlozEOSWrZ27n3Jo+8i8sNyBt0wQV35zm3OnodYIpNHmqI2hbvaNB/kZ6YliIpi
c9Uf/xux+YVypmfxGRd6Dm0TF1X3tHp426WiyGiCfSzGoqL7m2VckvGC0rlv+CPmKPeRtklN79IH
kdCitxMelCM1J3Oe4p3nwKc+UVckR+/zIenZplRkzd7oUkIkUbERtErr6FSlubVS+CgrjS5vWr3H
Bjx/Wfh4qznnrvI7gzZk2B8AerI7lA35iVtYzwh4fTADt3t8iX5/6L4LJ8EwM2haRjOvRhPjKVF7
Kq5/JNVRD4gXno/o8sZisRfi6ZADGA2gdCE+BEFWJ8ytX2iMzEk7j/Daw5Tk70F9kYR2dlyS2HfP
1VeBHlvpTxi/9gdcJQ02cymu7bbOOO9Tq5XaQwSa4S/hCuFDHdVInIO2eMywkYve2XGTeyFtASEM
1UGffPDm7GW+FK8zWBBOpyzI/VQRbiVBbnZdUAZGmQZvIY7X2Rc1OksW3QPRrIhehkQHqgHTEW2t
QtRZUBHGyF4gnthM1p2bzEPCA7ZAXfniQlI/Rc/oxFnYhw++RsEXeIPCNZozwJ1+RY9oUYBjHnja
xONCbm83WPQamKtdYKbmZKMgl/iCiJEp+yRxkvXWBV2jnl6THcUoRZlHwU3fyFm84xpUzuS+Q0DI
wfMdSO3xXHxF/XWFazhG9fHANo3j3kBffa7Cax+dB4PQA1cqrgW1cr2lud2J6A0Pjpc9GzNbtWrd
sTRjoirwfjVqatJkg7XSfpx2ZWCFPFpUpXy3zK314Up5DUcBL1RJ4V4xiww8x0xJ1/BoqK4+prrz
FDTNmuG8PhC9P4+7UkmF3vsckCLDIPMtVJZij73WhKqOX7MznDk6Ake+Ahe8PJSXIQqnY2Xmm7EF
H6WSQXHeuTMqsyar30vfQZCIztsvwqHQiXt7O6TkqHpwvqlUQVqJMaVJmyKpyyc48V7L+B+NnSu+
S41sGFRFe945fSl82XNPbtbucVcSG0yaBn1Bvo6lFxqudTYw2ZSYWawmnVrkWZrnK83gSERvgBHF
zi7klMRy6AMLsVpkhfEhsP2oD0vWachsWDeWA6u6NwqjEXtm1q7/pFAz5EwvjJBMD+CMXpRHFv5u
hjvy3PlkMN/OKTHT8nrAicyHSxRucm4Jl1c9PPBsRRDNLHu4OAElQJxaRCOipt2dua9cfVL5+tHQ
SHjUerQsaiDFEOxPopyfze9C9U6VMzW2jonjHikdvjm7CJ8a2EbRyFlqDWQnovGaUqcB9P/IVYkk
CdNYXvN4TylcnggFZvX2yHVYqA/AF0/oYzEyDjTJBKvJeF2pl+vESbqXtWE6oiXVy3nlv5wVUc+s
GUEtuUvNMUKNQQFccbDGgIvMwaUsnieIhPMjEkRE3zgj5HUs3kxsBizDGEUkg+lWu4QOhx/XoZ7a
rOtXWKPtfqTvE32f6I7zW4bF07ODb6dlUWiwrcLMF5ZTT4nYqtI5HhcM1VYtqbxrsjn+MTHuSBsC
OIGU161kU6fiJf22HtGztq+RvUlCvoK+8mCOpITjmxV74wUss8e6YSyQokyePz1uXlnWwQZsENnc
qMxEYm0tSE1ZcHeX6k0edQW7VmUxqnCTJGv6eetWVvLma7e6mE5yOARiQ93Tz7y4qEJ+cmWWWJRU
x3CmrX6fysnu243Hf0pm3yp/tjuVfcLtZtwXsB5z8PstUkXn6bwaZsiZJjoZ839FyFn0QusPTFGH
vDTT3a+WIVA2fMNSCNt5QUElCoaIUen5JisiOB3OsCycyoFHODcJO91Mp7Mvj3d3See9UpaXMClw
V6Oz1bNoNWXcCABfxbNEGzxay9ykts80p59SFj0RJT/7g2+Mxt1nJ83sfkKZvMRx5nL/7MXflqKV
9GpTek2jJIGu4LJSID9Ft8Km3If5dylDICqHCIN2/9T9s6gSZc5vgVSUw0rVccBJKEYsS/8aHMv1
WoR8wjlsKA14dN/H9hIwhX09opgW8AVyvD7fUY5O4ZZYUTi+Hv073nRMFgANkAt72MAL/JidjiTp
cnFHQCdrQcdBrVjirH38hYP0dGw4SKQlnFk6AN8Y/3weyuiN4thjh/wRB+bybCEQoGC6O0GG/xZ+
QLxNoE82PtlRqzYyZL0ppy8qzjftTnfn7n1U9W4W7+LPByzb1yAIKFU8tPQqYq14fIIRqbO5k0y2
+0i5RAaV5LSik3JDO58I6M6heoUw0VPe0QPRrCGgLC570ZAkwOMFBrpd/B1PfO63dUD58jWdQYV9
8dw+6J99jRQIMUg5q20ak9/A5U0Z8wBHdwArHpfoHtUPw9Ru08iFZTBHe5BtO0aTiCsr5ZeVZn1k
2dOj6S0AWzb8RXXTZ8Ybh/sp3kxP/cFmPbiu0H66f0G5mTKqw3XXF6d0Wp+Eqx6XTnt9t5fTZjbr
UYF8Rdfe2kJbnzDYE3HERFzaxtnIi6jBT3vTrXXmJOj6RUIU8bdpFNSm6unPPmg5ZOXpVcK8HWxE
Wxd+Si8lQHzlFZwQnOdM8iC7WK5RSHEghrqUsOB8amLmEL6z7vNuA2kaPKmntStTbPJwZazBYj7u
+JwsklwJzac/tgJqiJjKEUCILLYWDyn8kVXU6wG/3au38dwCHZ2cYNLR7Lf2KilmIKgdeA/mdOUb
t/kHa8SWWlYJx13LK3RUE2PQHHFle2eioCzJOnxkMMwkMwTUtXyQN8Zz8KUUJy1TIENcS4zby4x8
DCP/NS9nR/+Nh6Hxy9eL0uiaGxw6vZgO+t3OcWAGivnCP145oIw4g4OiAk+83LWGc2rGJQ8v8kaW
qAmMvc+9+/YDTFyaLPGFkmb4dBQJboMTtHEP9ixISSFXYZm6U8oTXTw+2tcS7tZ8bSffhrL0H9wv
rxy1TIIYWujWidmOclnEwV7Chnws54+tqKdVojdwnCeOOkQYwA+10GevW8beZUEAxKuoiV+1CDHT
CfpdIfwNsvhX9XM0CfeZ9GbyDkmkUsiA2cnTeAg864j800FrQcIv34rGS6sjMR7wviRz8Ks66fqk
qcRBtDTXP+lfAcZlM7xNTjszRvEgcUahbR8Z/xaareiLzYFhLgzrjSMT1DTiKWdIx8FF/IJ46IGA
2gLBPZxn3ETclL9QsVtv25ghJnueFLH30mOj56LXsRPh7yZ0o67aRf7FxcQDE15Rd8lGu2Y3AEkN
qkwskbYXidb8+V+c9wdI0AHnpW90moAFfVOgBe1RHhbP8Ec9wyqU+MsGOQHWH2wrhAxvBXZrfMe+
Ym/BiXOHxw83BjESi9pOX1BX+hJVR0tvOQO0VpVl/kz4cqD3/LnwSGp3XKPVfspuAWlmGZwG8Z5p
jHl/pcmLh4wWF57XnKOSXEIpNzq+j3hC/TT0sxyjb2hODoOqM0sDW7yjsXTeK/hprHVvNO85eMkh
zevUKlS20VlM6sUF2YUkjLFn9egWEuQ+mll0ZkL26IVMVUCq/VOUfwwgRnrnLkwQKpsucWAfb7W6
2/7FJEImPTcPTOIeFuUBqq2bNG2zkEJaT59SGqxgN9LNmA8WKmVwgF2yJLGueDovU8NMbjwp9oJU
Wny6m8KhKhgoZMpBW3njYiVUn8fgGpdcEW676o3C388y+PimRzPiiJUgv2eP/HcVB6+cbhSx4fJ0
KZILFi/vT1tXmamadmd9t758jSKPFtxCi0pfqk5bhHvo7wjPblSOatSF85TPeYQp90mDp5ivmvIW
KwS6r3Y41HybDUwbSat/9z4yOBLNZ4fzLjl2ZcOtLJESj0bHcP/0XCzoCAFWQ5Zuxq5wdoq9T9cM
65jji5zsVajtroWV+90JsW+Gdxv2N0pO7FuoEoIIYDWRSwq7E4Z21JBKwKLmfNcIZBNWooktcGvy
HK++mx03VGhGcrIE9MKK7MyxWIT8lSJHdyWLJ0tPpKR1ndRUQ7qZF9te8UQ1DqQB3VvIU5Uc6SI/
WdKPnX2T0TkyMjWwRJTLpCq6M+Yk5jzwVBkRNEbsJkkRGJtZEuaUiDpvstmTtn/V4Zv3+39o+Soi
oSMykh6npd8TVcYfrtJKkIxM9qJEDFauPQFGqT//uVjY6rZxchGy7/qmuOh3vbIiBKTRTvQGPuX4
8/OXkAHoCQg5zk/XFWB4H4iRESU4qGAU5RJB0Bqkz2CFlBzdOqeQbBwz7k8grUES3xbx66Adt91w
vbgQuwoOPiZqlXBhqVO71NjOd/3+guUp9NUSZw3MOytg0XzDLt/wSDSD6HaAmbyUCqP5W29DVbPE
KXU/jJjkN07audIBBO1WmO6cN4faQ9xOI50Q4r2Y5h0DiRtGFzeeuZNI69m0OHE+Rd6rznou3Ysu
Lpb/QOB7BzGsYhsLAOW8XY9rCohWXo8ugxyxGAyzshASLIpPeJrJ7fEcLez6vS8duB5vcHnMP1uv
79CEQ5k/I/MuAz+8FEXge2+Xg47h6MxkhY8ExFdMc2t7zRWHyoHW7WM18mM4weGw43S+DLqb4VOh
0ppInfdu/ntyrKSpno4A2cR8QdUdr1Tv8KNsvKhctRZMlG/v7JFb9AETA30qsSvP+nWAJIx5cLXW
0sl1oXGJMZmd4f+pZa5czMoFOLM8uBxhKi2ILfTiZX0d8hHhVJ3TMaP/7CKx4xO8QeImWqNedTsd
aPCoMrnSHbr3CuqIwMBjRCj9teTnpkcWtM+bV2glKJaEreUH2KIsNuiVXjUvwc3Vn/8wlLsyui8Z
i2jmMHDj13pXeDfHk/XW2r2JlcAG71YFcrQ9XJ8n7VxrJXCza9l9zxQIgevaNoKeGOpha67bl5E0
zYazz0aI4w6zIhllCE9gXFtx8ZVnuw8bH4e5bW6hgBlqww6fTUDfONEVmpF0dj7RxxzDtVcassmd
VW7c6L/SNvlKcKwMT4R5HmoTv/0FqKgvLbBKtftKCXe7KIG6TdvJrLOgCfim7bTT9WYpRLTSmB5I
ieX64rgGOytax/V62cCKH/0GxhIpU85cmgvGsPpZTSWS6eRXRLQB7kBXT3PS8PHpJFdATp1qNoEQ
y76Y2ggveyUvoubST6kjcN4hLv9mZiFpgh29506HQxnGwNd6CQU2xfLjcJCU/5r53h2IY+jfgGie
Eu/Wuj4jXyetEbB+DczMPrP3emAMlhtWIN62IyKbYPvuGd2xzHkbGb0R9fuSfP/0SU35NS4csTos
u8psqClzAtlrRFHEcwV3R+naHwhXxQTFUS7dSCw76Bc6AvtgtTgHGHOhiNAtynPjlZTZZvd+KNf1
hxKsDyrS1YSIRZbRVRp+HTlupekCiP5UVT/CeY6Z1UfsoiG2wlWPA+7v84AKo61mtZn9iF1BY1Ft
SwdB74Q1fNULbhgOZ6ADlMvKkd+A8u5iCsA9auOCBwmuN0YBNp0e9SAtQvzore4IzFsFhTiO3H6g
2W4e5vEoQVmcLlVm26QbS+A5cXPOA0wjYY8CW96+7ivDMlAYvqMSZ35j2uIix+RR0XPwiF8Jt48X
r+fZXF1rAtvAsKH1kY/GNpixNugEHC0uUxg6pxoEPCOJ175K1xQCI6beDmQM00nIAbdwaQGXZEw3
SKzCYNJGGxh4czRJLcA3H7Oi/gYrXihu2hZAQl+oaxtKerJaJ47Dc1Ic6OijO2LyJIPTjl2uJIjE
ru3xib+tR3lkOTao0XIsNHaHT9zcnHCo7yTPBJC6m+Rsfrg9+ZqyfuLSbIZJx/PUPD0bt8TeeXDz
QI5H6cxHbhaZs94JupmHxTMw6Mv60V+KWm8Lq6DlUxH1/HaghOp2Vn7CzPlK/uee07A2Xw6dq+4T
S4DPz+ZZ28bDYTOyKC984u0lWOjTSJOpCxH+VIX6uddg3eVe2kyrfd+KbUaXnL2JE0myiCCj/kZt
gTtcNGpibjjU6LcgIzj7pQRzU5btzonU1AlAROy6zuE0SKFoVJZXR0i6ia1xulUyPiQrLuP2ZaU7
1GNBaIon2jyOW0MNAZ9SmV1b7GFmbV9uuFhQcY8Wu6lu4utqYifwiPfuT6dTN7JzPjPjVfJHr4s6
l8v0DQbyzo0yPUgPWlV+sTj3mBjGWTtwgsfuHw97woq8lv/aWBZVSUClKWLIS/cvPkRT3CweRkc4
cMEXh6Tg0wBXK4gTumkYGAjiGWhn9OorJexJM10Cj5PiPJaucLteEJ4C0LwEHHbsZ2Fjai6ofZKK
fwf9gjl504dTIojIfXZrcofPngbHoMOhy2da12QqJKSfWp5Z82Tll7muHYxLnMYqqpPfnkHKFx/M
rRBnhbyh6gXyzjWtkE68jTYFocs3z2Fa5HjV8iLhJDOJ4OKa+XJx8SFptj0IOe+4zO/2CsID5/Bc
4g/Ajc47OkycJGwMjpYMQhar9gr6+eE5fHi5tbTqA1XstOH+4x8vqiG4PoaTpCbZ7HrW8wrHKf0L
SjknBo3q2W2EgpdF5qh/hx6VhrOqTQwSqYDI+Vhqm3cCjGetYnRHSl18RuypeaAK+jMhDqj2B+eV
NUHVr2eDezTvZNHxn/oCgKop5ALQ0Hi8eIys5/uhn0R+wFieI6Bj3c7CIlfyIaRgVcHVcYFOX8XS
KhZqcrMYnt4IVp3rrUXloH9YrFjbkfTlBmHQ5JxUTVSFDJHYyIeCtubsnIgRUYwCEO/KB/d09NYz
Nan6+3rNtgGZi1MPUo6ckMV806+3IPtzgqh9hlpD74YxxqDbGOGnEVNNGceKcKSCXuKLd//mtuHU
6O4343fAB22hHNB4fXWKijSkzmrIh0CbUGhwBYy4L9/w1REYddU+2ADfFZVjGvXrWdEnkfIwlRHs
cQmDIretBPELL065tDbwCHfQVZHxydkzzLrJcIIxvKMM/oyUDyE2e4PO6iH3OBwNdju4xuVZ1hRk
Ta+ZmNyMwEfsxKeVhZiA8ehHeD3Jw05XR0KM2V7TkeWq5UDF16yHNuVmGkS6XZyIvg+SnU0V80Bq
6iBq3MxMd1X6oGj5mAaVTp8+41Lj+YP8fe+Gi+VJ+O0LATueJAPsz+yC+k+C61L3fNor2PIJOkMX
GyrGSmfYcAhxoJ3OJwGNXCO1kaa/kZ2lbEwlgeR5NPcDF8c4wxEcyn8UBUByBmdGW+/cyWntjrio
w5HEuN23TVu5JwZH8fawWKYqQFyMZ1hYI0g0dlcHvv/ZAHhM2xfDzJHBEaVtX/80t21Hpx4Ug0FH
lHzCHuxVRs3Jy6KEoioiYeahzGe/VwzlGNgv4PFpLTgkPHw88AEjEDF0XDzK6LsRveWyjCiWHHuo
2QXBYqp60XqtXXJnjUiFutil2QgrHpIm3Qz6Wp1TfWb90JkqHEx3oGJy8795OpbOEzAkg0QJn+zP
XPVuZAiSve4yg5kKHgVabNUkiuKBAprehO+7Ryqm7SG1o2shjIxLCAfj4Y77ZOZywqvtjYwaRkHH
/iimlNS2AKiPkoDJJhM2S72bC5OdX/CUk1uuGDRxsCfKHUY84OmHUzzZRdnUw0dMrFWAVcAUlEw+
Dp0nvKhcyjBT/RaB9fsxQDZtTBiCkDlAzi69h+Yb7MOzD3dkoqPPmfKLg09fD9CiIvlnrP4yN5Q8
1Q6uwJi1FDr9mcH1OTlznlcz11B+sZWUgol+edJtUUGO+7TGqmzGQA9dipTsz46YRu1uqUKSk/k5
pDLOA9XQXkUwjIRYlPfciBfK67Kb72ntThfnTUqRU29I+bZzert07qa1/Nx5kE+0iPRouKyRzoXR
35xruN5SXX61TwGC+rpD+Asy/mGJ5b/qq3MXbud83vTBvb2kgrcxUS8aq7mJ5bzzjvi7aY3GYyma
2XKo7CS8DNKNkLpdra7i2OGuo7lLn1DzGoSACIiwbBs1U35Lz+ArgjppDROweZjmQqc94q9hz5Xh
SQOdQTXWioEP3NaOun4yg9Dw2EnWPg4VPPPvJ+1N9tNSRY9Mp5wTrrhAkW+1CKPEO8XcGT7fXF4g
xdrraJ9OWidHvuUzS0RMR83AQsIbODhuzimLQPSbkwdeTTE4+CWtgHIs0bv5VTin5UlP6mqLB9nZ
nSBVPLAYaYnUv6Gwz8ui/3xscpMo2KShfrNEcCciWBUAlSPAs9WS2yiX+tsmfizhxLnv+6ay4u2m
iJhWoetAriGF37QXIZCp4AWJ/ATSODsVQuPZgFt1M45Fabg084zwmq4zQzytQwQzuKelwJf/31cx
K9318ynZ1Uf+ZDuft7FAB6SjevldeHCjKzVr/xzJxRjVyvoUngMGuuhb2yMEAZe4LBAVWQCMxr/J
3pU+3d3lycBr7YSDvoLRdtYtxmJzKQCVaHJVvZQcH5d5ZZO+Km2yKqZaHPzVxm6aXIC+GxWBcI5C
gM5FmbiZ84CizgQPMB/i2n8maI/6N+vphZ4GsAw7OSe68UAoAmBi1XkoFY2dezY+zO28NE2YLwW9
45Rwir5buZ6Bh5mnvC50mVGkGeXTl4ykuoUnMUMZE2ZmG9pGLK8qi3/gRYlwUL4Ws3V9A30qc8Q7
rwUy4ASaufhDPrg5q+9FJ6AtjbJQCjAabK5OzaDPg1eAdDBP/zlWu4fCXuWaPznymPoz27UDHxOF
k2AMN+iM+y2/OlvZEmKFef1MYTqVyfiwiiJHym+S4+lQuX4Eew0Bk9MkydWHCovwQUTdPlOH6/CR
oOeFoxJZTxjx9N8QaFpq+JcpSJUMpbS3CiA0jS8Byd/udIShzsNeX/bBVk8RyYsUo/RGCeMNU8m9
mbeJOdFvGyUxG723b0tFBjUNN/OLYFlKlugd08/OgEbFsb4CYKq+vo1yHzcE7O+dugNhv9DJioSQ
NqTz+MIRZRz+RovUh3c2O3LDrhK7ECQdG/rG8wswIJMPx0XMHKnLe/hUBfs/5uZTOL8Gt0Rj/Ab3
UmYlp3KaqlTPi6MK3KaXuwoOqh3GH9J93hwICTmezeljH+p8P9hme7fLWi/hf2Hj24tuyry0Z0XS
GnMr/Z47mp3PgPDzuPtr10byjBUUF4r9jaUnm2L0XGt5uf7nNXvl2nEUNQSFRtjGLhqU7LrXUxQB
1KakiClbTQvkK0gqXT/iss47m06PATgQ0o3fwXtS3Dze5cazNfuMgZqwGHkpyjJoyblIpd0nIs4d
3MJRhYnD5I0WwhsWAMr973RZgjXNI2wUDkHnbY37AmCIIafJOPF7sFttm8+fISVcdVeg8zviFLwE
S5CU/B6rv3lpe2K9W14AmK7CrBa16Fuc/n1Pc80NRrmv8WexD4+9IFCrvaeP+keAQuwXL32YXlIf
kjDwlx0QvOuWGO69M4r6va2SipgD1hED3Y0Zc/dSFmBd1HyzzGDDdSFRRitefeuqJRSu0upD1kbh
A5giXDG5xoMPkW64lmsPl1Tk2evio19rvhwnB5g3MMqoVGwSbcU0mVyoTccuswmexo9KxOQPGy1Z
Ao0WtT5+HcIrVZlrvH9joARKRhq84mndvn+lfqwtiJHDXDPKG9edPcYRo8odFWhGWe+Gre4sxKLe
wjOCN1U8Xj9s7xpwb+Tu1HWTDF1o5oQDuqKzRYERUNhe8qJvrJYQqyIyb9jERV1e929x/TCEANL0
9cO/TPYON+JDBuUC4eJ2vF+KlBkMAcr1kOqfqb082Vierk1LuocP+J2Sua0V84vdg11WnBufGYSV
WE5/04/QXF8mBbYMh+hZ2oQIvn4Zw4BYhEaYBw12o4sfWpMs8JDlNzY63RXvd4fn/c01um8tNfQ6
CEXXIs06smgYaqKXnbZALr0ItAQ3T769IBK1wVtG5BPvqCwAioWJWcW0GNk4e1rHZR4TNsxfvlJq
8HXX4N0F/iiLdObVNH+N5RWhwQzEfLen3WCGWY/usgr+H4kTHPAo4ma5ofHoIZMasCtPGlPWKMFZ
QecgrjBNdMHLKcCIUcrxWam4zqLMSZmYZkTxKgItyP8FgRp/ZENza1POPFdYeLbjUhTs0eXW0MJ8
5n0LjYibDZxgCTYuChuloFF7lsCy1rGpkOu6ZmuZMb1xWlxgZDzRxWhCoZs5+F1PcG7aFyrszOEK
jc08/ikFTJenhTdtNA1W3CojZEdAFNmbNOTT58xu6ViABP+hWsQj9UuzSjlLEXC+VJiwQhMosij0
M2bT8KaF04+SVBTCKFia4swnjORPp2YQd+WvZPbzrRcWdt8m72mh74J/cumtIcCGLoPQlkjG5Pph
sIjk8EDMUfymsB+ksKUTuMte0J2bvvOKNh+W6RNY82YTAQ4VeXrbBuHflV/MbOh2l2yPIv+IGQew
Pqe28WvZpk+Pz0z/k2nxbw/Ecp0Zg9r72zoixIGXhsvhOGtT2fleSXN+MGVAppVddeZQI8kdwJq3
7d6eA5ZjzxFay9vOdJYy1KHjeRudIBtc3kO71fBJigA7/Z47HTQQiXf9cbyulEdHDircjpXGC/6H
njjOESiCkV5xtnkBLN5iGT5Sh4jTdJPCUT4AK8ad56gJoal4VXyoiPXGLgwd0zQwP1I6y/OQgPDV
LbtN6sTOc0bg1gzeXvMQMXb5QSA8fzrEltMXsSxJaTNHHofe+aDDXsWSDw2PWOTSTIONDszawCFl
Ia6Llf3Wi5WpJtL8ge/DKewJrvaoTDFuZuPdba6mRdIDXRPVHe5qdg+ZVtI9TSLDcNjr59ZKyEHA
Tov1bOJe8s7SOqsZZYRNonc66tJ+Z4vZtFcEG9Tpe4SachSfhHBRub0bQLapj/EKvw/Zf62g1IOw
nQX4qswP7OsQOZB/AZlcilWKf9moKWNWy8LwDilzqZ2nDqnfA6VTu9MMtpQXV4rfH8XEriL+Evej
jayG2w4Uf8nrgS9Z39IRy/xVTajrWPgCZT2cUnw0WxySrIjppM9nt/p9dQ7QW8DeQw92F0fCuQB5
o0wKXf71OcyTd6++CE0o/XC3ihMiYclsE3uhZan+K2oyn78t4hRH8zb5uwuqF9C8jTBchtqMoiUx
5dlDYQSzyhgcpuqVZgY/ZtLvPJD8KoBaRMMVYe87m+QbyLpLCuC/sZHvUvtWBEawbS2Qg1ixdbXn
o8iCx4sqO1yKY8YBfTqOjehQF30mhLA8No7qzELIjt6OS1xXQxVrH2nI3WaJRNcILpydTgYtUcR5
2bO8iSXf1dkBg5XiOtxNDf3W/cjOFaL0l4sRH+9IAmi0ejCv5YtO9HKSo8qrh4MtDQyJfxfcEFkX
cBDyGze3zmZynsHNLQIKaH9mw1ahQbtZK21Dk4wn+3CYB2lstkr05ONikum9vLN4E8eEHsISEmNn
AoLLt4aOsb6IelGk9kFty4LMHHvkvzJSkiuWkn/46t+gD3qF6+c61A/ewWhReV4Vmn9Lk2F6MwyN
ORLV0FvBzwp7uq7cQn3jDpzkTSM0L4QUvl7rO3J4ThzAvLSYCaVguYm3KXwwVYY4X36AAU/5y0K5
XiU0gXKk3aaM/uU6bNuvh5kr1UeEbs442cdFUEkHX8mzs2DZU6LEV4BDE1Qws6ccTF4jqp5lQZFt
PrwMFuvsob/Wi1Ssac43Ln0dTNjVAjBOaaJn7a9hdjlBMraMyY3GBl1ognfnHzO96eXCQW934gwS
LbpL7gQhJcjedbCipEj5xXg5Sf0M/ExWBf4F7giYOfIcVoppQ0LM3/PJsu92b38ep6O8RKpN238O
1fWrqJ86lkhPYyHZHw1YywFEdmL5fcFWhFnLn5BzmWevS/EIGJXSwHV4/plpuAjV3q3pPPNfmyQj
IVBDT0OGvVqoOU7ySSP/m6p9x5uApUs9TzYfvFqip3fI7E1+XOqY1TA95g6Uh3eDxPCVHqNGy8Gp
e/VI2zF6ZV6M6teaEhXWw8FJWHSkErCQEpXR9uwA2pNqRKFUhBRb21Lre9u+PUypZcDVGfPheOOf
vukKSALIHspIBGiMiGDv63fHE1M7DL26jQYeVOayGgEaGfHGy7zEQqdu17s9j/w2PM0PNF5CR5cK
3EzIdGsc29O5/wPjo9+QwIycfPjYKTXchHQ/ABWFtOc3W50rQmDyLwYJAliS6Zn1CFHFoPWeTaaz
sL5XgbMtTFiYABZZcESuOqXc9s/Yu+uzWwJSmb+NX/sO1ujPpcxJh3ZSccwokG9K6E9FJ7hQqZQ9
Pc8Gp/38PBdWoSAN3h4APj7dN9GLivCdIFFcUO8yaNwjCWexQyzYWznlnf4vNqXIirET6wYaV1/c
prCFcDNxclWnlIlYrEwssvPb+bIMr+KO7oXjxDhImqwudXfvljaqpI8L/y34DHHgaWkJGTOqO7AI
f7Jwc3fjg4lVPCdTq6KiczuShtMCcLJMwBNsR252db1HbontSwW9SxRihLfRMbw8pU8M+rwpzuzl
SIeAGUcySZMbDd8ee6t2Du7h5aTkNAKDcuF3O3nL+6kjXho29sDKXpZuyLOYdyMgufuvwiit/A0C
L9JR29B3z5FsbZieAaNg+/sfggEGgcuakCHtfsiFB54JMTmoYrdZ+3lpYKPeLku5d1JVlzShKl+i
yubnSl11Zm6nDIDKZ20nlmTrUc9Zsf8oWAH/BKwed/t1LqMEcECo01Z4EX+s5VqFQDKlc4ZNEl+E
+gVKj72PP+2HJzpoTNvOGtc00ZfnK4iaDelvVh+2MAo0k10WrU2vSDaf7XAaJNspGNB+MIYThhHR
1nZLkKxDmKGJROD0Ftf7/snQlfHZWseCJJyzh4doSkDRn4q6l5xVIDZ69fR3NkJmwF5E+AA8kfRX
QXZajMMDvg53WHOeOLeilU/9zPUt7R/pe03grE/sZpxzPFiVZ6OO0Wj9Z+WKuMQhgt/4LUobU9hz
NVzh9GdzvY2YJuJPa9K92A9GXIEIxgnDS+XCj7RpuQzJdyMyLIt8Cn8NHGtTGSyjjH1ZIiwtHrjm
aw5oK+pKyY5c3c/89fxvqcflmm5PYoHN0UflaseqTqM0bqZ3ggtGLZeBz7BQztF4lnLiaRa5epdH
J7eRaydGQE+dqmpd9AtbRF6s2yojl9KuegvaL+BKgJQWGQW8H+n71uDfBYR5PQNVGY+RwSDoV+bl
qigixH4btebZGr5W0AhcKnxigiDPZa2lzBUBIp5H0AoqiQS9RtVnI+62rhZqUTcPRWmATmXMyUmF
zS9T2c4jPYp9UWB+kduPvhLBTsdunDICPAU7M3+f29A1JiAT5bTwnbgjoOhWKso5dmfbzoxOiq9i
n8/z/iw2O/81YP+T8TvBzhUZOVR8DH6ALkM9dSYYlvOz1uLSCYLabv5PlYAqMFzB/ravxBKir0Z9
DpwS9cRI9l9A8zHKKUNLVa1NHwUB4/WIDvUROisWBXsvA1qceMZGNea6Ndl1g5TRTirklDJdemYl
cLRqLCRzX3y26W9c52jmApFA7n8FdKErWPblhXxiaOUtev4OrGimfPrDPt6FxCndGfFL/uZjdnAY
RSb4O2QPPipPTIT/SZkyqOVVQsyg5EYWv15cRfmsNTcCKwUTz9H7lY86VKqEm+KPVzUZEpaxLTCN
4X7SxHo1P6DQnIwXBZO+3TN2R790kLNYYOQu8MQ4blxMQ5Xkmc4IJm2X184HlZHsSZ3crPC6TZCG
QwEFoaBPI4q33Ubxfmm3gbDIwKR4eNE+FnJhuJk8cuLPbz4MZo2IM2TAdz3Axz9W8vrI1IZFRNDF
6zg2H3oiwgJ67Fki1834QLvMqcoOYHHyopHy75kTciaMzXdJVpX3tpZtWAhzQHOcy8EPUupsNeMK
N14Bx1SyM2S7TMFX3IwSjiOxyv4LEkk8MAmaeyKX6VP49bZYoR7Whbb/6vLKi3gL94kvUi+BknLI
V5JA0ArSRU1T0cRdpngO7kXAgVZM36jYiE6F1NXiYlzHnaReG8l5le6eCtOSSbrZcrBr2jy0DBem
suN9UEfixeQhUEYhLNz71MriWFED7cpZcTkOFdGPJ7UIDGNZPl36p4cl9XWGofU3xC/ZAmEhf/no
t0D8fAOc/sjsMVro6tedSxWvlbwHESq6x5A7/TafnME2t8eGKOLpR3ZijXbxiragKFqAbq3C/xCc
cH6glhcKF9jBbzL2qf0JRcIWvgHorqdSxsiHjM9YmXm+CKq+jo51ngltg63frnyrwfY6i12oztGR
1opsLTmjfX4yblG3Z2xNn53XWUa9xJeVibEvzow/lnIewEHHmr5H8mu+EaC9DVr10g2VCDWm00WX
h08OuMzTnFXLK0nI+DNFZyHtejLNtMu7lz6Qqdi4yxTKhUAbHs/3gsc8OXrYRTtxtOPzuQeDrnzJ
knHvfDi6euvbaoWj4QXMvhbzUVGCG+ztxkAJwfyLF3N+9BnWv03LoBvy2VZbLaKZWNMbKPpcWRHO
DCplKorc/PJX8YvJ96fThW4eL7sBEZNWY/bEHv0Lm1HWlTKbLlQfmvmTqpgFkwtSkG8QU4Q0zVHJ
okZKtIEWtlRdHDcc/5fhcQc6HQew1AxM8efSWMg/Pz9cScsoVKQuLCaz11xoDC0uAialOCeA/NY8
e1QRIVvyQnOYuP1Zpqro7X/bwucujA7NdAsblVV7LSWUUAes+gcnWSdVRRgoKmBUEPPdnC2gKue3
lB0/wnfSM9Z34BkfAOid9Yc/XxM8b7e/uwnMnropGR7MbUB0SKMYwBq/bhWCdPzpSPGUcWknkIeO
zAoAa1QkOpyOOzD5hFA0nAqPU7MqKmLld6GReVgb+URg+6AsjaWDwgeQ9GxeuvHGbBKMAokem/++
d02UZ5r9R/qK7GKGT71IeKQ0LNnAjjkrW6fgqelHjMvORmddVXmv2lp3P73ZNQOykD3uM0vRtKoC
jbBWKgrpUG0iq3QMjNOGAhKzyBTqt2QmNyoGSWAmhfW0NKwbZen2f8J+U6mAIssBnLp2+wpoklNe
0uUKa+jzL7UL5P7oMjq+KhLlMkgk6dZ8lvswLnrxjZedeSxZb75bjOpLCAyhMk3aSVXAkhj5bQ8z
f7vzGyUwu2/AEzz3c+hQJaA6lLWtWxzfhKu1gOIT1ouHumZO50+mKhNsHhC6XpsDpDYo0MIJ9hJy
Gh3x46Q+N9Jkoqci08+RUcGLLj81UctMFiZe+cB1E/gINxBuj83jKisMzoK2mkbU/r1vTlApaHsQ
cE2EeSTMDaQZMuFD8NNu4YDI9phThuqiRibbhKuiGNbPXu52QJKuohuXUI1kz/1qDJiNsPf7IGV9
3PInUl7y1EuAPP7a1bTP3VM3ulgnOB/TaARxxKJejz5sAZrm0HaC1D2y+qIixjd+kdyPnKot0Faf
abmEf4skVoU9ntAjiQyhPaRSarTmF9f0ppaT+U7AwtKaF9KqdV5YNcBhqJR/s51B3zEQJY8O4R1f
YUyq4Ixxmi617vobCprIM84gdfDCv8ogsocx38ARagoo9EQQ5bFv6w27Rxw6y7U/oXf4PfyeF+Z0
0tG51e9u1ucecQZUEln8+NX/9STPXsoxoJPj3QL89MXebnlSYp7H8ihYrsYaFWDe+YK1gj2T2BzB
6KsW0eHTpCgUMbulDbKlChn/WFZCkRpMMO4jucP/HAY5J2pz0SU2mkRiWvIG6UaFMZHy477kDxph
XUkuprncN+UycRWGmv+uTdxZQ4qmzLPWIF4wXHqoBn3n0fZy9ALeIemQJoGijacmAJY5dDq81mkf
vgQ4gxQZlQYYqsZv7yLSRxsdnIRpwXBPHb2FNGqkXnQyZ7Lpl2z2GSdZ5JHgTX9HdxhfgeJkUSvh
fUkrWHQB3rHFxuoGinUnEA5GLdDkfKCS+UEoSweCcWLyYdjCSzdzW2KaO5Sra19WGnv/bz/pTmkf
S3K2YGdjOmLOFh9yap/CW9I4ysKU9jpQu3/Paeaw7naLMCmew4LqTTmIcTdCzBsmuoXXB3VaPs3w
aqv3a1eTqT5/mlhwF1kqOVPYVVT5mDFcln4iHNNqnjrGquz7jrEp0yar+UB3SvXS/GaZhxUiuwWy
WTUy+cdC2bB1JvFEqYQ/HfNwiQaScb0ybbKwv86m7CbGZvw4tWYU3b9DwgstTIZgrCW+hOJrVGSq
kW+QeNseb4jUi3vrC5ybMrDic+iahDo39fzAICVOlwqGQ3fVD0kZPeyvMKK+MSbiHQuRkOC3r3Di
zzc6Ngb0tqo9YzBivG00yopnEq/1w+JHho5cQYj5eRu6oHUR/2hntVhneF2BD4eo3X130db6SMV/
xjizA6ImbNkaOtD5qUUCGmWqaUzU6INlDWXcT8T8MRkNgpT48UXvrUtsmsBfCvosIuwTMprhbrCK
BSYqHzaIVGfLKlojr+uXTVs4nI9OyF3ZIdhNkYajr1eRyRqjLWrA4m5UPKRrFubaNxjlEJanTSnd
nVAFI1B3uACP8tkrmRLLQMa8avEOohn6+NndWzT6mafn/kPL0JBh/zjqhM+FCFa2xNUu0rW0+klS
HdMtqf3sUNJUFJDEPMWLggMpBSZ/57C9DW4JwHNK6/F81+yMsTAcpTjYu9qZCOQHseaQ/R5neY4A
2aQMuC5CVg6ryWRHChD4Hw2oVCmkjb7G4FotFEXo/NcO8XD+Nglv6a5DbP32QmghSLUjZfvZS+kO
WRUY9G5NVbQgyUzwO0fF9iLnfpzlTzTuw9n6utZBlupYkx/2wgzp+BKwfZYCic+UieQAQB0/z3IM
LYpYCMhrTxkonpka15qhqWsmqBQUkO8oIZeLkQg02wzGyw3EhkM1Grh1mBXEeZxO89UhxQI7ce7q
w6oDr2W04K1zK/xKSJ0/jwGo0jLObZFdqnuO8NVED6xgeoIlxSMkV8EjZunS2S9XATmc13Pm0e8F
7n5plJEH02uAzTXQ+oJ32L3ZPf7tcyMXQBejbHVUlya4RmjhRBM1iYplO/cbLKKU2DTZSHuR+4Gv
X/b30FlC+iFiWzhEDcSxJzHmFO1WgweuDZQtzr1w1LVJmejUftz1DzdUePQ6oUloEqmn6voZWBeW
FzarwhWOcjw4O1S9FZqlYXJV2BS0S4QgZFH5w5h4sMNtvjAn+GodiExestBvIA2KXoRuTNIgUeqz
KHV6mJGXEXTFg9fhVix+qL40jzxWYtUNJogO/n39h9Rx/oYTsWSMIyaEHLNzWYYOF1H3C2HIz4gR
eSOpB0R9gb+3I3lCGkUoqxwXb1JS6eiyz3nv0SuAtC5uc6Hh+4JlK6NGQ3LRbk5HYoc7Vh0incR6
hihOTCycxBn6HfRaCU95rodi2TRN4ri8FBLriafcOt6+4ZTojwkUzsknlDONu2K85FXOyd4fCvXD
HMrJFzlEXaDGyPxyPY+GQpdp2a0Grm+Mgr0M0le0OR19dy3Dbcr8EfQNttuhG4rmr9aisWZPilv7
bRV4UKhzBKgfGSqQKaSbvKpwAUInQPq6+MYWZHWKlpJY38i0kk40hcrcv4O3jjgRpE+1QLssa/oD
7HfQOjA9SQF87cw62+9+QlLOxbFwkk6Rky418P14cd+ALsdN3KJjv2FMoq38FKgr8PLkfSDPHbmL
6ciNEwMVMn1Dz+v2xxcFkLHKuTqVHJN2po2T4LuwZftGFXgC7t/cJb1faUe95FWSABcMCRkZFCk+
daQuv01042ezwQWoyu6+gZxViIR1wR/IqlUneIhFbToUGPSEbdZz1dqBNaC1RWpiG9qUJsU0phE5
S2IotIc0kTVpPDuPIoMOzUUPm2zmJzLVfWGp7JCYzJad51rG3m67A0IlPO79ubtewu4zvlm12iXd
IrpoZToa5pvuqH5eUNe9raBQHZWqBoMwAXvx8lRYoxsh5urVlUNZzTjUF6fpQxoWkL/KMht1G6tr
zpDImYx1YXSX8wZjTA59LObXDVdMzQqzlUAPvv+MOn24x1pUjC+6FLo6+IKUaxfStj+W+CKO4lQk
kHxOV8dRxLlu0irwMPcdauXQheudJzwoJsUqF3S8VgIyyYjdnHeN09MRHiVtra9i4bGg8oNhSec+
0ic3+TGJ5fb8PjjkZIiqlFkoMEU7jFJ9zWRREusWJgSYpkWUIH4OFUGrX0ynefgteBp5BXxdtzse
6cdNqvQIgCVcAki0c4K3RO+XJrjNcF6G7AowVJw25xN1pKCprMNlcxBE9MCU/G/lhdSoo4pErrTv
OFSb5CDr01u5nE0GVkzggjOtrvX+PAjL6FCCuzuVmK20sjhs+R0Q+DqnkiyFKK7vuS6Xedap/3oR
bii4UrjmyWmzt7smt90MnLt/FTQPKHEGKo8brdj14ov+1IHakvuwWnkbQ3LrDpSY+iNdrM8Ri9nW
3+CJ5NO95j9pladr1GF3G6cmoI5uVdKDsCZ/nZqnc6AFdzhpjzOYdIXVhvoFXtk7rdtt6qlOLwPg
5W08EHZPb1HdxVfzUU0y/nKy0O0LjICeOKviM+XTzO1oOZ/Nop1OZpwomwIYfLjGDChb1T/gU2QI
iwPUIMEALrUmUek0vx5ZNdh5VIXmcSb3NknScYifWi29HPu5rvAKl3QkUas1m2ljjJpC9ak2p1Q6
UK4aAXBu1rXGbGDIyLMfRqd8CP8SYzTjjM9U6YYwWBaQYuoZysl+KmH9I+tag6WA568rab2JMIbq
1vnjnAmY8DH1DNtOqpXx8PQaMJ+KY2timXOqXdJk7qrIRKJz+AlGVMfomEX6nZp+f0XcZP6ZyfEL
Ih056cIVOuCGnrlDjjIcWUAAhylHQwx8CeAnlEW8M5CHhiEQWlAc/lW3kDAP44SLe+LdUz3q32h8
RV/WcLJuN9NX98Yn5oSh8MOGQYCJdeyTsoeX8cdOYwLxXZzV1U32BkPMaQw8m0Nl29Gh0GIeH8um
ue+0DQaIbbXSML0A9rHzXLYUYNxJLl1Dgd+pc7AMKqnZfWNcy7VVF4SgfO1Zj5g8RQGKaruRb4gk
21fT+pb4g7O8HAjxY1s+uzylyRhUJ8sTnKYRb3rFRU6arPOcFYkLl3ry02IgKYQ95V43NXiLHqtO
6rT85kYanjWz8LGcREdDsjGvyLV0aEhMJV93lj6oTkM0AvlTkqRVZ1W+emar2sFJXYfIe61RrKUO
/DOkwjh8Ju9c4PO4VFjcq1bkvY1PMi8PegaB9ZiITA/xxFGmB6f1xzwB7oCC6c4u0QSS+G4a+mup
eLivQ13+ttIKvUbr0G/13j36ofrtN2mYoo4tQy8c4GrVW3MlsWPS8Mwz5EAXfOSCbYNz6bV1j+uS
wct4FdqSlbrJT49snrdl3HjTHu7u4BO9eKsBt1SeOCCUK/bfS15cCLqMjKAvSzJsvXu9vnKlTtl7
RhGeBxhmGF12go9M5Qh66xHxes+Y9KlCD81RJ0MVbmbePHv9dH41VY/zXio7phpbAUE8En4lX6+W
M+6glLnKGGEc29yTjA6NQGf3R3h/osfyoaYZmxBDh7w/l2tazs+rPtOLCP968v9dw4TX1mvUsp8f
DxhQ5frVz9Re0szLe92B8F6UE9933Ae9Hdd12YCFbLPWPsTKG2o5LTr7FZ5AyCM2NTEnSj3DrHlc
HrJlCph81S8dGWdUjckrb2aj56ub3p8bupbTNdNwRx9yiOeEF67c8gPVc3u4PbCRWoEZqJlTPYl0
e8Lt2hQ8jU8+QFg2uB1Ei80447I5VUW1+5MId8Ppg4Tz89kNp6m4mJ64fKke9L/TX3ym+ePu+GJd
fnJ4cWP69v+iBWqJwMrIUwsLZhNTU5XMEjIsncQspEmXbWF2CqsJ4h4ykwc91X5kyAF3DfofECE4
4mpcPma0keX9cSSWox9KolL7FW8oQ3ew6v8urcON3Z/HPBb+n4ed2zaL0SfL/tM9Xd2gaSAsI2i1
vy7VAXeGFIWzglNSiymeLbVqe8CaTnhiJwnx0C6iCyImwx/lE+xGCdSnVXzjFcN8FAwCaYAHBdz8
gQ7himReEDyQWjIgpe0X2XcwoqjgH0+vzHvCmuxO9aycRn5jDNMWUuQfamc04sM9K1bGIldMsKnh
NwC7tue7MVZ9NUua+mxZReJINIVXCLbdQky7pzICcL6cj3HbD2vvJwuG/I1N36DaMIte/HQukk49
GX3gNCGHxo8RAwI+h78EdsGlkfbfg1PG9FCA+hulzgAmKNxX43+LgtgSX7IB0WAIFPlVJ9K4QLTP
hIfbaJXeHqeGlo+ZumDVJaqp2erry8kFFG7M9lR/RJiO7SI6+Ri2+uGg2lXAWtk0WCmQoOWYDeh/
vxJLPAo09WjrMm7LtHaGkhbG9kNDnOIfRsPcspHWB6TfFWvyAo+F30l5AZQ1Pb4MJ1Xwc2VKDijm
rNX9vaBMJBEwgRXrv9ysVlg1XOmEP4kFR579j+kT9DOyNBQ1hWtD++u5o/5WsS+3oumGolOMIilJ
kKnssbQR1O0nxL4DiG8tlucrorjo7lCqkLVZN4xFy19vgPvuGxKZTVZrcQ81AR2cN4BVB5Rv6jsa
Az3XBWE9PfbgrAIlhdjjNJLxz0IJkhJLtE371+z1rsiWSvjgotl+xZnthoQMCGebnp5ga9rTZwQB
VL3LhlKGCHOQJJsEf/5/4K956/MQBzEr3sWFY27fakU19pZJ6zCV1xNH5ln7p+K0PfkNQQG4ynTp
3+SPiBXeXVOJQiA0TnQB1lzx19WupVKEq79TrItfVFKTqNODCJLt0X9Q5tWn4FOntYhMMn7F9W/a
aoBfQkJjozZzk/I3BAEhWlsksH8i8dPvs801lua/lR3JOFiB0jtS6vYRa6LOWPVdIFKLf8Gg8Ak7
Cp0xLA9NT3cAouWrrFxLpr1Zjh5xxY2a/bYYtcuLgt1Qn3LtGXanopmWgR7Mky8J+jU1TIhEeu3e
9dbm8k7xMR+oSmmiS8MnraxFJta6Hz5jL0BKHkukH3mA1l1vgjbf3+KhRCITq0EsZPhwX9s0wW38
R3IuOd18KeoXnX3h8xzQJQ6y29tf1YhWs+yT3bvvME3/jplNchB+sw2FgQqEjbzWkd2SuHJqneHe
kIBVTjN+o2brfC748ekGfCLk/0ESFPb1ptuKh7UG/WaqlfSn6qE3SyY/QVurqQ0lkMulFwI6LTPG
wHtIHXXggdx0XNSdJe4xzCn3EpAnvQB8oeKtHdK+lLIa2QMeszFn4d432PR24unc9b84Whxaffa4
WdwCauYxaCzVVsAETVolWV//GD93rXqLyMw4nkIhur2edp90fXi77EwEDt1gobwhpyZxNB2lYmrN
XdildVPzbDkUwZqb8oez2+Pk5YoXMTFQYrhlwPicunvgaPJ648MObBCy/DMjCgv1Vzs8L/5u04mu
1Ns49RA2ym+SN8rx7mYfvkz2XrvEHPSqj+XUb9LOzug1o8aOEr/cS1Fssx/PZfFZykyfLGMoo9++
goIWMMnySwrxez6zsypwYVqT/uvkhm3Swk74mdgkQV088NwPWKKM++lXNQk8n3+e3wnObsJmHkSb
GMBMYZzw9e4Knzhms9lRlH3UuMbV96Hwhh0UokJajalGpkPcd0g7xnhFfmRqWmKsl5BKWQy92p5e
xS8xev42mJjGud4kLLaj1BuBKqivdA6ttPCN7LNoI1MMAQxgx0LTLyMoXJFiRhSMeGvXRR4iPy/4
mEh+A2nHrNPe57srTT7P1N6SfMP3DJ1F+FCkl9YVsjlby8804gT4EBTkbCI3dUrv2Z7vu/nwxzOA
/h9efEWwbJKzszstUjwYj1hFSlToXNFPX7zO29dvA6Qo63UJUrrV++C7e39Db10ZGDYJmmOkypRF
ZLxc3MYmnXPywFWnd39Rfb2sa24B17P/EDy0vYGYanVoP9Pi7Aq/U3R4jSkfPxtl+tQtObNciSIK
eauho/4JE9doqSMo/uE3TiZLwSY32JQxulG1SEa5lb33kX9pdIL6av7NNmNKbDtrTFcsYGL+ANEP
vluRBcfwgYcHRnRdxMTVALQol/XfDdRC8VnGsFMnAr7M+QtBGAb9bMFsz9ra3aK83tTEnxNnkotB
o17O4DWjVM5drQwdJkSsO+NDH0CJQ4TNmIzqTKoLB3Q5hk+Xh6sgce6OKQZN2VOLMc6cNKOfv73Q
b1BElJlAnfI6IfpMsDfUIMzJINCn33aMB6z7C0jj1fnzPD7quearWAO61i7MCpY32Hn4I6zUGsbz
m7OpLEJUE3TwY1oGg9oY5RCX3zsE5jmd9Zzg7D7dvxXjROkHrMLZtBphhMJ67R1UZNyKvclIacNl
mBlfMjXzb7FGR55/g/YVYeZva9WWi8zD9XCHQ1HYEEOk7F3D4KImiWyA/77W27DzjRMHIMd3a4gu
EGP9PLlSDDkSj53y7kkJFPht8/CTfDaEvyFn9UBpyPM3hT4pIiAKo2/Ck99qFI0o6LI4dFWJZya+
asU8EJyMTD/4AgDHg/nmTEniLU/TYqJs7YtJ+ZLMJPETA+FBou+CI+QqvAoSTTY4qjEqo5hRb1I+
J2S3OPlMEEs7JKpItYEljxpKZH1BeJ7nnE5iM8/NQMyy2IMy/vmeypnnqgXKgpnJ5s9HWAoyQRbF
bldlHUTiCcLsXQRSqj3CX2rb4t8rHCTFezbqVO2dg0iXfoRngPgAxkGHZH0+58jGV6Y8lPAvo0KA
Zfr1uEoctfkdeP/T1lGXRgsrGaFlZVWSAxPf2XjL0CBt3AeGYa8aorebWQco+hGx8VE3BvLYh7zI
x6BzEapxV1Fi7y34xF7AqxxdDZHkCJLI94+hNwNgof+cC6PwtdtLQHWDHJIcLW7kHoeNvG3WL1Fy
jZzXTuxpOea7cgnaUyVYt8JAjgieJDC3jTkae/7/DqUrwS6f9G6AtoJ78i0PeUyAvJd2RHNhgONJ
sJJFjNCj7WoQUHZt24uBm5PrmnPRkailyA2jsWgJGng5a7jgqE9JbYBu/pfF6EsxBBI/4o10Bjoq
g23FgMbrVlrKI3LMyHaz3BTzlmrIZidKDYFpwqYhbOMAgxGFEEktp4PeuI8VA5/ceTYe087iOyKO
Xch1fqEES2Tu1cfjpnlkfPCbZNmxzbJPsTyhx1IOcwj+pydPNbPboiWObcLKgB04FV5FbIUA8Whc
Zcaix6+H8clG611k+a+Q1V+d2zC8x1UtmRtT7oetoQRG2DUAOQhLLzu1cKtRxKQ6iCwBdRaq0Dhr
ptoYdeB7zdOKrWttNssFXYLlBGNx7b2R19IyyNCHRTEin16LmuE8oEHd5oFHxgcEIIz/kiMxsr8d
9JI036/xU+DCRY9mPyFUdfzQMOLL4Jpiq5bc1PPWDyDQfDJAz+enPgOlomQsjMcgjRcjsWfyMRvq
3S1W6q7XQrB/LONwKSd7LX8gVom8R7jAm5IbL7FZSbVRqXC/Duz81zQ3flDl+lNgKD5h8o+f3PRY
rJslYOPk60GAt/mg0C8H95VtZ3+2HjtPI99KFiZCp3H3bRl/QGjW7sunNtJfJO92RYFUIUVItLPk
9vNCqNYnphSvjZvfoXuWUyy2fZp4t5lnJgU1KbiWzhka4kVvPR3932BkYjvsUbHWowk59K16501g
JJ3/IotC+sz8kTbqAO+8ltO4WgSFsZk4ThdV5syET8frDfRK4AyG3rVqGs5/6PgUMbBdTceGZLv6
ZctOX+pdUrsdksbjf64jGoTcR6AHZ7A5Oj4aeZsdEMzu9i/niYrggZY+bDaxYWRJjzEktOTd6xAr
nXNs0veEMoAYC22EQXAE6vJVGIuv3KQhVsB+YnXKSGU5U/YHOZov5nfAmQNUUDXiKKQAfaX8JQHU
0adJWbxWyk775/VGJSzDqTktuZDf/kaDTe3WvNaXTMHJcUyaj9bNgUce+YaqA67DW52GI6TsdAos
ESciwwdgoRQM+uvRuofKtqkQEOnkgcVEWC9WaVI83bdeFSh08Z5tJ4SNjZWF/FcjWgvgZU+uhHSh
+FHR0xgycHCCorMbANnp+R/ruYmkds26lFumZdXhYBdgDJuQt9RFbiI4XLLEDL79OCqcSDTBcbzp
0JByHN2Tayiq7kspenFGfk7muSgqY/J5ZqpSOBM+GNeS1XEXY0mMbHUtJa9yuf+IyzLrPwnGWfkM
/QGY271B3kE21O9AgNsMFb/DnabfM4N/tQbHn7pd4E7N7hy8GbXyNZFwCGBmP3dPpMsSHTWOzDzA
cswa2StjFn1bDC7WQVj4gthyE2Xk/WO2KYlXoDbMq+k0sMfdTpZjdmOYl/iX/yp9BlVQg6rYmyAM
eRYVZKGngND6Fc9Y3XgRR9hCQ90b8jZzIwEpc6Dd93U+hdF+cZTW05gOl4L5EwYYZRA/Cxy9S1fs
Tb4gswmYW7U/209vh5hbs1MM74g7d6GoQjwKyEeqWN0VL+G25whC9AgBCuZW7O89ZLvDRVmk5bTC
fOAXGHXJ2ndPERcJaFrzEaUP7y1xT1qXR/j+COIbZtn1mjIpQIHMVG/19Wl5fdv+Zd27dOpbV/XG
/DbTAQ66jw7EEwHg8N9PCcZjVAsfShY37jrhsNKK9nfqPF840Nphvz5fQLOqCGTA9eUF1MAzy0Hq
hbxOJ6HkFqDSGBVUv/DovMsvixsdSb4vJyZehcJMu3NdIfTnK69UJpQ1z21zzy41D9P0Iux77LVq
q4+PlKDg3zkdXFrZqqI2shHGhbEZ+i0I0JPVEIb0BNOyU6iytkL/yL/683mTGOy3jH6+/Jdbtwdi
YdGJh2S6lOd+DK/BFny4X+OG2qa8KFnzaSbKSHBISmsRt0x3YvgCH5qu14QX1me+WCFEQeNU33Z5
Lv1bj4djZbgspFFzL3RCqE27nK5uS4ZYWCOX/hYqS8us79PkAQ2sR5IquSvO7ujmc51dAY8ul0tu
UFthaz0xpTDGypNMVRtHN1DRVj0WsKJmb1YngqQNzEnLWhm0iu050p+ahPcBow3tnzuOAO/9eKG3
TVMkSEZWr66PbyqpHoXkLbIQ1sK3qrsHM9WTdVxnW11phZWmZvUw5i2BLbHeZaGrRpH1fxPQpbMU
UjECOw1Nur/4ZxNl3Afr7+grLeKrXljdwYi54yYz/uh/lWu9os5ZnBoLRnwJah0YGKr0gCXyb6G1
AkKw2aiOgxYpJwRo9zBuOQxbJ6TizbOi9VZhVfNPPhdsb5eILdSslQKwmdHDjQWmC21GrsUqyrXH
b82O5WRUVLUOP7s8RM/13TjpK8REc9FO2KkFVeuw5/60QI1qlmWfK8XlTSgCJiXDuWaoo3j7tJYC
hsSfyULmPpK2DQBDXjF0qmS2337aNZiXQDKYDQmKKBfiKjI+F9PFBuHpVBIz9GinQ93AuyKoopN1
O6sh8imqkmeEjn/gJh991aujkRiEV6FG3DFwR4D4BmockcSNGIInghYnGeP3KcqX5QBZgem7y8bG
dgoF9oQAlPgt55/nKu2dUP5e1ZGkaTlOuz/bdoi9lwQ7Ryn0xCYkc4taTE4ThVptXRhimguY2P94
bskKy1NsQkveScZsHZmyHuMlFxgs0lG0UeHArIIw8N2vEU6DDCBbHHGt/qrt28Mkcv/bpsdGe4Hq
6pAhf5zQ0MXkeNt45acH6cwqaCixK3sUdJwszvGyiRBtcGC3l00n5SY9vTM62GPhHPGiKp2KXRDu
dN+MMu4ayytRMBUdM9rXM2NGqoLgibI+p/tUmx3CmGNn5dix2eIhimPYBF5kw1Q0JA0419Iahhtw
XiWGBzaNSoY5PaYK4GCQFrXdQmTq5CTD6K8a1CWMydJbFERGzQ50sg86UDuPMGd1771vhWzQ+FTX
wXkKeAWlhtqP/+TpaPSa4nIJCT73TD3VbkQEMSg4QOIFFy0IdUr72mCG4ycZmAHcBVOC8K9wilpP
DIlEZq0+M8A2ocGIpiEwhzjA45vIgvPEVOACs0eZK67oYHlbVYsPJDrTrky2CKQ0IiSUpOV+IiDI
Zut8jVEfxom1DQea+tGTmy3P83zytd5aH2EzBzOIqlVoe6DKqml1IIBtgLW8nSQ9o5o0RhY/Fv0o
lPtDvT2ENS2IoJBGAg3ZltlpBtOIDToEBfOHFMbdrIK20Gq615Zy4UUP+3OvrZL+fR29KGdFbaGL
Qmki4n9bdvMMjdzSpNfwYuk+ilW2LpTCDNz/0WR69WexImRs4iSWnjziNntAY6nWpM4xpl8ckMq5
8Fvjq4CbQjI7hdJosQLq1/6VdDONNeeiIylkK6Ch0QQ0IKMGD+LU1cBCavgDyetkqB3+dwxaxSsO
24FqdGgVphxhsNaNlNvI5JkkCu9J+FIDO18g99+xLYf0aZYFOHSR8XNWsuvyELxfhMmvZicGcCTo
5JeFRzByjZiypYmqWUigdoHM/JWBUkFPaxg3O+HFKYxUcOmLDdDAMPOKfxbIc9iSVJw5Jisqlnvk
6sz9JHRF0GsnNrcLZu3QTq68OonDpsQ/Q97H5GlUQFasxDEDkaIqqr1fYkE5bYl4ZUsxxdKJGmYq
q0UrDBKkOyxoHnZXsHCYU7Uy9dW558YS8fgnKfzSGx47/F8co3RtHu2+tpAombvv7oazQO6dNNCS
MX8GgrOp0lYez2eECy2XumO/KbFyUopc6zONYZoLw0Le3LzCK8eVXs2hSleYsLVGjgAuft0Ln7mI
e7vHay0OtQ120ecf7UXrKenaO73dATxR14Yh6tWCqNicIBOe5NccuwZni+nsZqui1eCGfuRyTId2
jDba/ZKPorADqgC5CUJAToMSh0lMfGHzNj/in1wLao3h4TJHf5A2o0GPwqYplO9CyjE/dAVkwIgL
diKNDQmlS7Wx2D4A7UCWOL54uHglkA9ZPsgVpDUiUJ6XQcGEKWD1VFuI8eYZsStrIFwbljVpZRZE
s4IKGfY63SAMMrlxWFr4jczDuWSUIBzTzCFFl4IBUtuER3IZ4yWWdfNf4AMA30iH0uiyNbOGqmRh
Ri/6t7893CWjBDAI9Qratazf06MkT2ZwXw1xwUIP5UzaozV/aXcoe92z7gjlK3zqgJiGAxanxQys
MuyVFqc+arB1jWxWORzbWptgAr40DedfGtlzujKhFE9z9sIZigw7W3HdyeKOaHoYkBfABGOi44om
zrZ3aQYjQ2kSgtahfzj+9cgpOMV5eu66RWIepvbbEN08lFq9fcbqJCjwpxfLPw1vVLNQ5mG9zIFw
J9bB4qn48Gg/m4hk9A/O3iIKEAOyBLRjE1vQzJjHNrPXfNDUzxlEQQ5SOrhOtVzq/xPaCf+czlBe
QHOMXle7NWFILBNNJoY56Hc8chFfR6oV42S1AnfgTc24HICHbv08eUH6d3UFQDINdaj4s3rzEb55
sK9qRSd+IXyKfk09EmKkBRVvr5PMiKoJMaT2He2hLAoWzF6tlHY+4aLc9DaE4WQo+6ViMrzYznkC
fqpkmaXQMDCpXdNdHGhWPhwvsnGGBmnSXVk/bCZTpQ5IthEzETGY0M7HpDzkeDhM6GVLKd/tRzvH
w5EN12qJKkfo9vdwfqEHCoOQlXqukGjFooZZjnXN3wuaIt/k+QRIS+jBVQsrUwQ0B/VOZckw2wyq
4xa0vmkn6eqHgFNwl7+rB8zSrQ+J2NzsYF+n1vQ+UdNeAlfjfB3HmP20jeUfCLTemSddLuHXzQ7V
208dzhOeiP3bFh6+vJWPimmqG2XaQFpNt7Z5IVnSiWnHp4gtFc+SA7WfnrUOPRcliLOYYkHQRzYK
oIVPrikEeBXOMia463rkxfSZneepehsqYJOQTiauxKsildRZ5JTEz5DyjQVkkkI7gMRQhgbmVECy
3h8b1q3J5NTfx21WLZLHviIz75Nfccsyw5zl+TOKWNRUPlJTG/2A0R4AjLEfC8RexsJ6ts1k7PG9
TctxuYxsrn9LmWIaDAIRFZFig2BirysRC2Et6xp38YWEKwHpBFDtwWOvbGgos8YLG5rDKJPH/xQO
hdfGdJ+2QbV2Mc8CdzaRDHtaqPwq+p+CgwSqz4urNw+QNWshSNv/Cdvf20fYFfY8abPZKIDM/YWw
4NjUd01O1w9UC1SMcH+8UsSeYuIU4jkHiHRtAXqIBLrLIMUHL4Zqpg3JY9ERzmen2g9fRI2DSSKn
jgEuMCdVtigmH5pLhejcFV71mc+i+bGrjwYm0Y9crsc1dLDdkAIpIy+dmkG5fuNZPFa1XCMySirk
iQmqdOnNK8xpJysQjPCEz8PSWuGYmnt5oT/2vG2D0j9ROoW54Lk9+RHfiqDoU9jqVrYgsLiKI4jU
gAklWHQOM1rFdZaQ/OL0VGW5mlM2GOS05cIQyxjq6CoySFr7FQraPKxTw0Vw2JtMwKwjQUzXy33t
iHBuNoXq6/FSxZdZWjwvLY9TcNrDo6tWj2pJFavHA6zv+aRrL/Czojiur4EQKWpGeIHPBs435xWd
+bm+qpruQJghKLZbt8RCfh2LU3eiBBsc9QLz3+HRy/0fqONSHF5cba6UAL/2+2+Luxo5sdE628I1
YpVQc+t+PpNvsYPpJWjN5cOe3qArw537yAi9pPBC5OH+e2+RsqJaPFLEKNLb89XKt+g+chjeTVXU
VnaSdVk3tvPlxM6f7/RrLyqOxHxkNrT8iOpHhWyuvpRfd9YW1wo9F2QTByOed48OMkGsTbZ3hI9o
ouzINut7hopNhyelSP6YECg32d7CZljPhiZaxKm5srmC+cMNNSdr/8UjB/lI9eQ7uWIRZo5GWfTw
i1RNzSfHudNVcSqffgBBF6HZJA/wf/MK3tD8Tb/BYnZf7meZlyxCf6ND3Mg2Wbvj9Tdxt+gHEalg
mUOm06XcypqGkmyM1MsK3Q+pdQ21f7YjoPjfTokbWnPkJ0gfqu9ONTKLcN7/YsoOCOPsjCHB5DGJ
k9yDi1XLdPNKZKBhcS3w5dPLHFUfphk3cQopxklgFlkQCqQhcR5z2DHAmAS6a89b+wBIEYPvJVMg
g7N0BSKLTX34jq4JkvujayQF1oQOlbS3geUM02K3qUGR3HQNjtLJpOCCMWZFPbvvZtJ/IR7pxKoS
OPC1+3/8QN5iDDUtSH29GJ1tPfjl21IA6jYPUg416VffuCTbnjssagJg7BpVXvjHoJOjHCuqqXFR
wsOhPKF04cVMcoTdxDnhb9I6LeeiNiEABF7IhLHJJya6ZBd/0OsT0pxS6SNpowsTLymqd4Txj1Sa
3UBrRfGO6/M54+t/5p4qcYAAwKJOBmm2NNw10EgV4Or+AgNozG5d4t+KTSFkWdLl9Qz0mD2pOYkq
wAvqG91c2CiLxP5OxrZLW0tfSCc8BmC1JahZRKzatv2CzJx63jVSWIcPLr8ip1IhEGgUpjEbwz7k
UAMOlQrtwS7jCT+0XwWYwl1mUa9vxrp8xLmXcmAGQYKeIBWzfZh8ZQExEcX+00Pz+LDWrhe/MEMp
l63z9umGFHQQgtHoo1ZuS8UpYxPmnpTh86hgdScLjj2rhLrTt46fXhLgbwPhaE/NKQsT7DJnaFvl
rXbuVHcWW5JUH844rj2lLasjkFGfJqIHN+V68ys4C7DC99SaPtuOJugAgOqUO+UNzj9Wi95G4uBc
0SgU4tSlvKKNwKFybwMaROwMZOSIlhsI3D0oOsdPpcGThVYZdGtcFHlbsfZ2BAfrEo0jnwyniKFv
Lns+PlOuCW2/QycIPD0os64KKDA5inDuq/ceSR8xzmD3Y6aihrwMjC3w2Wyr0yhpO6E2b5hLB7Rm
JjlBFBZfVCd7Ys0SRSN4CbkpM8AkMOQm+1SbXt9oXQFk/XH5EzzCosLekRMZmYjNwFKqMb8B3ZKE
El5oEPStUfr0V5iuU4QK2UovsswBafsds+Hs1u9J7m67/T1+x8+l3PSmXALVZbSOupVfWpVct/Vi
K1DObqBNS+BTnyhvnBaSvyG/e5borSAIpdjHKrKaQkTrCOgv2W7BhRwa6ZahxKoD+fJQWq4HfetK
eeyFKSHuEHYUNZGsOUD52at3+fIMY4YKb4AChxyb6Flr1bbrWECRW+r6qHLkgAsjrbh2t4O5ymiV
6MG+8NfBcQ1DqMIVXRUsQxsOQ2MmMPOd8UmJUUbTNMO/8sO5xsgp5bEnQhy+mBGhyx00CAhmvlsO
RUHINnr1wvCEDmgwCgpIGPucP4rwhbmnMeTxOdKiIR2YQq0z81S+MbYDkcrhd7I5R8gsTJsB+qhz
7cfKfVNpHKGU8oZwBwTyyE0irfDaseqdctNMsut463Erqkz5mfK5ESxaGB+2yfbGMTTWh3gHAdpt
KsEvWw8iLNV5bWYG267PQz48nlJhX9jhVMjmiXghASxW/HlIkND+g6U/wBJosStoREXn6dKUx8Hc
yOgAQjZb6TjzdW2klKxEViP9m3UjX1gLNmrwCTdmSnZkN0N0nxiEcLVBOoWwCPajICrxBloFisxm
wccqvAgZk+42L+jfWTrRWb1BkJ0dJmyGXerAuhGm+gpq6g7txMh/7SFMLNFe+aoIVbWQTAkKZdsB
vw3fEsPZtF/faHKapQcF7MhDmUCejINOQrdcsuQFzAejHW+Q9qV6KAv5z8CYGKxm+3YvTl+yF10p
pseW/tjkf0Z6Se0GUg6q9GsOfovuOww2Z4Sb6eZvBWJYOVsRfzeocpIowysjhsCW8wLVcKd9qlP6
a9EmOgfUhuqYanwOmiWK5cS5g17MnLvbfiuPYM7L02AEMZo5iyeWp/9YG12IL8XVOOQuIJGeu8Jd
zHqk4ux/WqD7FUXiLbpgeWEAFD5qBVhaAhIzG3ngstLCxPdFwn3uE/ii037HNzDCVA7schPkRylI
x8mo0GlrjYpaUdt4kvGxz44XQc72hQrDo6isc5+wRQGXo6cqI8n7fNQD1fIz2fMrZEKH1oZfn7OG
D6DfFs7ZHjfhMR4n35BW66x8uF2Gdpz5vC8q6NB9lFNUVFjxCuj/HTZA8gl3BUPEC+e2J3VcEuB5
9a3b3GpzhybgwD6HbkKL5jYBJU0CnZqx8xMH2/vcBVWYLRacuG4jLYS8eg/4drz14N+7ultxUa1u
uUk4AmN2O+ubDBgTnAxDP13Vx1jjqJDUgsSgkqAMT5+rjTeIzoGn4aei359BlQ8FQ2cHlYa/03Qb
2AiRsOc+MnBJvOUnq/AjAVPIQ3Dd4jSDwK+tdt0tpLurKyZp3EmseIuXI+UQHm/BEPVxqFAm1DCG
WIL0npSAH2/lN3ubb2yWiuJZL0G5DBj5eWm0DGoWwFaIb3HPetvNf0RUeFSmT6nzUlfwKYe4wBrA
R2MTX1dH8TESDo4/MRFZ9sSI/qsXhCx5ycs0sSijoTT44ilKj6MLySMX6WNhqojNR9bvphf4EH3x
z8+aXk1z4sPJMxdUX87O/uo0GI/Z5giboMwbiMbaUy6MwNKOeKjtOG03tUNMgRgAaTeLpvmOf6nk
s10+Mc94kBdfUjnyEv3onWONaI4PkLfyVn9Cj2Nqh3w6fXnFwlSwEx3TnsFw+mWjooTYChHnE8yX
ip46aSczrd/GGLJsnmkwskoLkAkbp+0IPzea0RItY1RxGOjlRd5kpfNpMBZHqP+zp1SiFss5VCdX
0gWfvI5Xu2y8TG3zMc7liZI8l55vCtJvr44kJ82AWGHqmzncGhatC8abzJ4utjtlwNSx2+fTUFAQ
U8WAOHe1NJXwPMGrVE7DK2JDrtYuIjCN5zMwGu7BzJk8bFacx7B72ualdKan0ZYwGfktJ/osc+ve
pJvgu2bvUfRU8oe4a5ovltHSYST77e4ba0cUa51S/bzV+8bQ3ZJORw5sgWoC83XiaNLvmx7lpedc
fldwBtpK87KfV3xuMlcc3JFuAOCgRBeUZ8blrnOps8fQsSUC4ZbEH6NNotfVMzdPOyu9vYXkFz6x
3UrPJ5ZxoR3WWjgKhMxaL7D0/vjsni4J/zRua0R4FD+y6kixPQJPrhH2b2asa3QOdyvRvvlupJXs
+7tWYFwG/y5U20xix0Q2pE25cjTYifOKax7q6ZbHxMbtRdoZMS+T3xZ+htwQRqmaYVvA2jGK2inT
BJTcpJYHeYhOLM1S/O7WlZat9sj65WeanmbsMSETcPcoeIQ6Xks/SZummEcDa1mwNsFiYVG+lSbD
n2uqdEq7gC33KznEjXnp8JpcmuwzMbhn73dVZVjaWdeLHg7E6ccWMg1XDpXxOlFiNIEzMG8Vopjc
EN0HnAY6hXtlf8Y686TKbDcLwEaVNE7SBH74ccHCyLAXP5WW/VI3QQHYANXyTXiJiq7+oaW6NurH
pL6UP+GYYHD8fslL9ArtJHK9ecbnrwA8Jf4p9b2gWoYTh5WEjR8ngICDKnhLRzT1fIvYLE5PNZM2
NdbeVPOtWrbecJdMwCMyB88duFo5gkl22BekIq8L/iPQBQc4U9O22282BjUS128LiVsw+T60rGVE
yoxIv7jMUuyfHGn2jQV5Lep0oD2RA0eOiaji3+YDeAL6pEh4MtLM0TrCIVF+IHcEdAqS0e2ADkb4
aHPN7+bF9fxBxCh1IeoSj73JZWKR/oHQtt5cWPBwMbOehOwvluQgZ0XMn4LtSI8hhdms1U2DiPs0
TwR0Hy08iuT64riudUaiZ4J41ghGgvJHK0T7SfjZAd2uZFAPWr+lGO9dy/Zd/7Gh2ae4VniqFb5s
FuO+onfC87Ge/ySaIiQwmAwCDnr1fL2XMSVO8ieiOWAadQGL7IFmta+0H7ogydXCcK5KHYQplIWU
f19NlOg6CE4ji2tfovAc/k7LLMitG13amEc6reJmjdS8m7uvCF+/A7GRr7jzGNzixTy0nQZ07L5Z
MbHPNpwpV7TiHFeUwmbmkMeGR0PVj4U0zrgnMTK5T6gCYgFqedUkSvYSkokPHEidSuWmjPoFn0RW
SQHNXpo/ScuGJkPIPJGuDipzlf4mymMToHUZLMjvRPYWUyvH+la0m/rWZNEaugM74Doo0Tc0zljK
CIlv1uxKwLVJaqAZLGOX/e5fnpj5yZ+hpjhVEYL58DwYNNX7t39FGuXY8BJgQz5XvNo1PBjR/cbg
yw6Sa4CVtrZWIIBEFJXKCQLcLZziJI/xOV9j0xfAkHE+sB+YD7j2IAnG3Yca5YiKRwtKZyhpICsL
PhSGrs9XyS84G58XoHhf3yVxKKejBKdzxhi5qtADYcQ0A4yKLX9X0bM+D5IkCgXz3+i4+F4Ng/cS
du6fULaNyFqch8tWlnIbdk8xTeYhXAjaee2Yo7pbZIwuZKEitDcQmPgP3LxB8HXpTwqIM/msFkX6
y4FRX6E4vcRbxAifLOjt5rMzzvpbqMJPyEO23CZb66bRGHYGCu9SI707RnI4LmBf7oeC7n5u/3ew
D3nK3MWSlZ86w07Vaz7F8JBzA+5//9zIjes3OUeIN9/E7fdczLBowBuKZri80DprBLrCjitXqNTQ
noyFu/QHgKlITfFgMybIabxd0VWnwXIIkIG66GjPapX/+lfDA0msrySvBi+T6u8Uas04FmF+TOcD
rNy/WMVFBuZnfg6nKaXRFN+//KkPiOcsy7NqIST+e+/2YoK6ZpdcQ6KhutW6bHuQY2W9tLrkq5y/
DWKJoYUav65VtpVf4oG3B1efiW11SGpdLoy68E0s6aR2T0L72tS53xpv6++7Moy11wlcMM0BLTTd
BvbcqDGnFFxnvFjYa2RfMiiQYXncxk+0toNCRPJGgH3XyhjWjDpYR7ofr+uhomv4gy1wfxcxVw2Z
4Htf6KkJsy5+m/6rRtKUYcl/cDgGbZ7f3FlP9tY1cNi614MudpmQvFBNOAciceyLFQQFGmFMJ5fw
ysYA8XgGTuboYtuCQuY68J5hLmvkb4LQ4cIoQcz+CuKlmd+ebE7T6UuKySt1CebMfhnZIPx0t6re
2Sjl6rZ2LsqOEWWETJjP2iqbzmkjdsEYf/HqlkpDHY+bn7vRqgjNBjqZONz8y6+zisqvZ1I9yfHe
rLYSkQ9HZVqQzrHImsWEy1kA0zZXHMYPpTQEoVYNp9vMSOqrcB4VUvNh6mb/UyKcHxgDDneg4xZb
K9WYqAvT7HpPxKIEMj1u5kDXdXZ/upq3sL9xzvxLk+/tnR+2WqlcdR2JQae77LDGmbbpmjLh5pur
Ov62L6ahAR6aLqLibQJWCJVEUp6uq+nb3CO6E34moHhLD4jit+a/Qh42vJT5AENilXgLyTI7hKjS
5MpZuR5uPmDNduFFBwV0j4F6aFSavYp2YgDFk2vFiKCsQXSqRvygKXHdd60A23WerS9asH6EMggG
6nYS3d1xt0zq4XhOjl/HcL/duzf4tORzh7rLIauaIGEcuDUyuTdpDCF+Fu3VHA1Q9aZTn/ZloxEe
c7ZsRI+jWRp+refGACKr4lE6dPSpD5o25R4GEwlsio1EEsyqw93fsaFOMOmoRaf2GfBESx1ySXC6
PuhSArmBJpJx2YD8/IOrmmLcb9OBwt0bBeId9wWhYBdvGaFZhIgUeihAQdXtt5RJ+zyUl5L3IWd/
glDj81QQoNVPqW9zrQeartozxrpz9D9n6hIihO7UHx89DhyG5yLKSkkAcoQNYq0+H86AlvzV26cL
cCieN0NaVqimddDnp2c95nlsBU8ZPUIibQ/j9SduXWol65y4w0ZR1SzW5r8WjIIpJ9Du6vXWGyXN
5p7J/1EP/Rd/dydEoiSYIopJPUYqHWmeV9I2kwo1UQb8v13B9ZaQAzMf679l4i6DnblGnvaraiIh
pFfEEPS8JsyqsbTMrfMHM/S9WKabo3xEcvORyQ5B4tk4vB5v2uMjff6Ik9KfGeC/BylFczCIaMC7
3cVdMxcXpFPHjgKiGvXwZ/Ge0baGdVTcxzdMwaovkXEvyKR/YoFyUApLVxPYS9Bn/ypfiM7Yvbmr
4NBfjG4hXjNTrUJgu2AuQfxlmauWA7ckXbPLqYSvXQpqEgqheM4FTqC5dhUx/0pzUdwFxA3aq9Qo
mjrdZ5w8Cawn2AEgqv1uj8gBrBER7Hd1QpkeTAS5/sEkSA9SXB6NdtKmMl/PIlAJjlhu2ZVykCgd
1klWFBpcyR9+sXU997DDIDgvRWOLGVTnoCN6RL8rzttE78O9BLwZ6vsEaYOZ6QixItYojXvdE1Xo
WiVm4fI00vGAkY27GrG9hdwj7H37eW/Y80B36slL/YfMcgX94Gs7REyYLychzkTXv6ShUy+3XEeX
rgJjFIdDL72fR6MVGIpizfzG7NP1pTr9Nsn6sluueCQ7DgUnoZkhmihBQY7zUM5+RVOcN9jIuE8V
s7IfjBYi0bJNP5l30WNp3ecxb98YmewOfS4yol5AriB4eXMYz24Q79JOsXWctMz/P0zsNcb1TSH2
JrLaGTbLn3UM/HxHBOF7cVHtC/xbpdRd3+MRwMqDXyDjyIbLgkFH1UV0VVyGEBl7vPF3RmAQ8433
vkA7Yz5X33bxqIWtrSvmTSCwTVK3l56hcMTL6tuzMOGt5xIPrUhqY+5tnHmScgaoZcivSo4g6KGD
OFztHlXURbsw94m25mU4nHpp7g7c5yZyxcOM5WwKnObF5P12NAodz4Ot/5N+aOMkh5kJx7gkSTO/
e8wRNDMTvjRKTpOHLSFNPxjZ5KT/AlhpCKlc5Ox+33wXQU8xTq3lvHmzHaolI0fp+OO5Cl5YxtAQ
o2D00yJ/K2Qfse0OYw/x9tSdW2RFfCAdT2jQijtZxGQI/lEIbQjt3H/pDPv1vrAauCCruxPD1vdX
5YRdXO9FSL7GLtXUlsUDAil2/sXFXHZttNOBAGQMW7td5HsRTNfhHy2W+wnNh3JfpyAU3SA29qsY
+eMXWHyeq69tKAev3iX3jUfNS+twuRjcFNipwaBBMdxfpKEXwtngNcpLQ5/xZqxWdCjjySDHSqnD
GUgGL84nwof2XHCkO36IV7knply0RhP8Kc+oAv4NJ8Q6bjxPh6z8hm+HV4byQD0uWKA3g5ZEKcdD
SAsfdgvYqcqWMcHUZdWPh8/nB3ndFaPAMvH4Rz4Xq2PNHuEzKznKFBJyFMga6bBd38dYemb+XVYR
0XjWomp8MK+GxrSSMFOXj+KRlGFdDEjFPQ6XPmvGpaKbzD1+y5sMTZMZrztL7VsP+pCxNgIzVuqT
nR1d5ZQu685NsO1xinw3BrJ5wdeE8SWNX5EECEg4536MxtLtLpTocdzrnJECeiEOsU+ZICbYPQF1
U4tjrAYTgWHbSjKG2V7zUM0S7QDRIEoqrkRp7zuW4e+8hSExB/ZBoM9WAPsF3BIdx+It2pCj2zon
B6A6AYoU5jMPYm/m8h+cjyacakDZNzDXslBKjyNzMTGAfZIVtvTGnpuABzaE0P3M9KxJc+bkVCCH
30HUV6FwZQrURHDgMuc/BhuN3LT6WpfKUqoGGEuiKz7rRODFvEIN3MV9VMERzgBOspJhC7QLk4kG
OyUk8HwOLThx3FKfasjxpToMJ9bdfCuiwcAUPCGcMLUdhfeqpNh20F+UtvJGr3eJGm17yTI7ujqL
uCGGK2Nz671a5paUkZgu36RDh28gTzmChGXNslRuvpUvBD9NmCPRCQB3AhzSZyj4KRTFSOK/6BVP
Qm0LtimW2cPxgRj6FxVxG/PpFqWw4yxEFouP04xm5U5xDAQEqyvcZTUOAnJFLtx1/ZAT4M0C/M5F
bg2vHetBweclurYkKB68eHCIE3xenk5Kuu4jvt98/phoOn12BPn75rrd402ko+xzySnaG03oD+/e
57ummjlZbNX1puByIyij41fvIHPjsVE5Y+3CX5QnwVlPH1Jt184CBNTUfEUgROqhLUN+XnouHpcb
iYRDBttaKKQm2rbKqSbwN229BVS/Qd0rlOI4QYLNCx2oZVzzI45DuP5baHMSp8xkgPFKvcRQsdUA
t0ZocbkMnDbYJz+dalsE9rr4zKVnmgo1VEBQUdOS9mYnWemmD5v4GiS7rlCJTAk2+uNbwBJTF6gz
upWxLNh/0QnVnhVipuSydrbXzQ/DSf1/Mx+kZ4vDsP/82veqCSsudk5fiKNEr0oDkUXHfBC+69zi
ChTyN07wGqrALGrjBvlTLK8Duhn7PkcZvM3WU5h/O4hiAoR5jZrCfF1iKCHPHu6RUDOONk3ueuPI
68s+l0PK69XmbqQk4LK6hLqQf1SpD22ypKtfkEpuAOz0O8SYlJPjXdc0oFMEX9OoAIS63XNA0RLe
1q+++kPmcq0Wu6AIbHo99UcRuaFOkjXijbp/bs/qj02fNlkAYv/Bm7MdGj6DWgDi7osN2Dwmr35R
KsJGG6hNFVa+6x+xSRMHn8fXIWai0kMmEAdJTDMYj3NfP9ST31PR1zuLoGD1LJJJ1q2RNvuiCFUt
YwqWDQeyTqWuE9oRptPSEJ3UsTYI13xwP/Gqt/OHXi0+NwpEMZP1LSr0JQeQPDhR9+5C5LP8IpPp
jJ0VDZVYvk6VHwudH7n1k/CMdfnTLNWXVr4CNOEriZkCtFredp3SXG5TrG0loN4DHo/YcRZIQzUb
yvJiTLnOyigGEEK802Sh09ftDvTZWu5TulOZrX9xGjf26TWcH3rWQRBmZr+Tvk/VU4PbRd9m4lLq
sFfaAvblKjyfD2xRaEig8zZvHHS2S5hBmXJanl+TmBv7YqlsEvFSFKp+es/mwYYF6MEd7JOaz/WA
51GjyILOVjSx+NA18wbah2zrT4oOZ289vGgZzG7glTmcbKA99siZSup0ifyHDJVVp6WmTBqkP0A4
GZgr7XPD2mlCA4lFMwHJHIoezgLwdi6pWj7UsX77oqzXJktcEfY54h5TOH3f0Eb11SGFgLcn3VIt
SQhmwIHKmOybXtfZZTQkWxc8JbiADRUisn6HY695X5tS9TQAWoWPF8C5WNS9eagR7cKCPnlLsLE4
pnuItxB8R4zmXOpU2enSPgkX+5XIPzG47CbcjTfJM3mLdUyk0bFb12lBoOS7l4zjh84BDPjFq6x6
S1sL/here7UBNQNLlN/Pq8Jx2Tth9EBVf0/QvNYBKewp1vXN7ytMYwEDCxUl2/hFysG+acNOitZ6
f49nDX220QMC10+3PyypulgRUA97+H7FzouB5SfSKkYEvO9A9XarLFoCJB1yQyiNKtaMuXQG+mVm
x94GuWdr1Znzdr6K0XB29KhRnzsyQZQvitFhzS71sgfHaVj7VKDajJPeK5opiy6cwYJJpEP+yfl6
HhBxdxNO0SyBfVASRopuOr2TSC6BJopuICouQGX7gr7VOj1Be5hdaxi4vZdbV8dK0rSGAPviHLsJ
hCqRmrAT7WyDnV1MZUF+P6NCs4Zp7dlYcP7xNUjikonhFzOcbiElSb7CgkekdxuLK31pMbPzBv8O
a4PlN1Gi8HtX3mo1rjUOg/kP4O3lk+V4UVDw+2OqVz3M4WmG+PVOcxJ13XMZGumj13/2xkG4fdLz
zyovUV28MQdTY0siZElpCgvzWjxpWoJD3I+NoXkNUohue8To2aibrCjyTODP6uzKmsE1B+5LREuN
w2GT30qFtZR5vsXjjqfbhCuR+1ZZkmrgi1iH3RXwEQhfprGNMes0fQaMWjppPYPzGb2nYXH67ETn
F1LfnKnbkbjW8FB9E9kZ1Up/huiq792InpAUCVyECZ6dqUUGD2v8rgyj85ZEUQpxjWRJ0qk75MBM
5l+cJUE8ViGGY2rmEjGPkhevQ1zEA6cpkdl49S4MGaoNyM9iCVTBBw4A4+DuEATMFxvLe3oOpHJX
t5JSKi8aAJZ14X4OIO7RJQo3wkHQys9BpovsJAlfq87HoSspkjow1VW5LIi4mWFSVbcz2jTvguS8
kOiJh/IYIf36BWe4wq91NxjKSyVZFPrNApufFCNbnxEcJgEnaBpGgcWMvcyU9NXuxu6UdSmtdzpa
OiwMVzGyHeavjrDp1QCctn4Ft49CimNPUMN4oxfcvASJ4dJDYLtsujYzuUK6W3pxh0GNSiPy2oT+
yUstVnyzTtpkJ3om++FagR4FPP2nk/RNJ46+9Yy3Xmr4w8jYrHPpesEUKTV0fqPnPYfH54kFDqqG
V9qZMYdwNkgSR2/ZNDN/XSU0HEDuQrcRBrsmnEYoQYgOTC9gK8CBR6cM3q9/RHjS1kmzMqIfqdVR
k2tqHyUIzJ1sBucH5avpuUWM4f69jSpdRKc1uJrtkkOse4V8HdskvrdjdxblECia1JD8PjF8kZGA
K1bY/afJtslaEhkbaJZj8HHLGv8pErcUXDLYbCTIdPWuGeX4atJYGaDOMuQ7Hi7TgxiGKyLDpo2g
LZldsEa9oyDdiEYMhQwUXxxJutW9DqWZjB5ToodnNIx9M2/IOm/bm7FzvmCyCg6Q3Kswnf7m+rAe
h1S7D8xVhhopoCgpLU5foJ4tZ4R0Vc+ySwdveS/9HTN1CJLa7DJTddn1A2qnK2zphsNNwnwI8zqL
qSTPLIJnEhJRfXdnSlAwRI3UmG+wFw5gTXJ2/GGyef2RVtq4llerT7QlpZNa185NONpDafqqRbk+
EHOHz8b541UKf+PTAhuaoM8SZXxm78pmna4MC0j3jaJRftiPyaFTj4jhk+mthPGZmQDpEnupLBLf
WLf4Ty6npoSef2bT8ca9EGDBf3Zsd+y0zEIqkQ/DJfNuQr3OaE68LkmHcty7HZPWkKPWuOEZDN04
oP6IWlBBanQMRDdVfi4c2YZ5FvzGY/gagMYfIIRrqzyz46XcB0c/2W0yL8Ppgq+4bGWM/KendfIq
wsGsvS+8HbcCv28v6EjTOyZ/aTmzgtBm0iLjqQ6qXHNCxXCKcpT/2S/QlZrZivgRhjT3qLnsMe6b
+mxbyyww+g5oeIOiNZnV8c5R53A53Nby8FPwMLXRYn5CNxYWcx4GrMaxj1/hxxIpBn0wjsyLw32z
ZmFMgTYeqDhUfLWDVdK1YZv8HFSNl+UDfHcXhvQ3Soaa3dppKVpX+MpHkFJSO+GaXqRpnWNuT3W2
ydNM6qcOB3XG3Fy5ijMcKqDmqoGSKswqmlm8HyDg7bdKbvWNjgEidd3OMWFfhWHc0/KAWMyWdmHX
OEM1XFy2S6y6ICSlD9IF4XSynmjAJWFhV3x36FkFarNmJt9nI5eg7cUOoVsv25ZbOS5UlToNqIPX
+w5VU8uWYzCjfOoFlUxI+9HS/p7UKESkX3wbyFEqVqSCvgaB+Iz13jllJOBYLtQEXH8IpLcyIviP
pKYgrj5K+qgt6Iq/W8HcXfuSuIiuNxNq2KGiyoXgr2qHJtVbCYVFaljAgfCxofuABEGlDVP4ftMq
Ou1pZ/8bw2FaiBpfLq8bjNwT8UUrttw2ELJVxizUX4uyGGNNfNItZBJ5u1eVdhoCUeOCySXegCMV
Vn9yDbIGWYrH08d/hFM/vJmabiGk4HBEYFrAAB6xijcys7tCpB1yhTDtCrZc2vfGhh/A1OXgAuur
nOGSM71Dv0D9enR3BI0hBKpw1atCoJFB50kHe7O7fpL+GZfOAg+Q0syJEFyZwZj2cFPu6VHFUnne
jRb6TrKZ00EmO+n6V9XQxi4kPAJ+IBOLoR9C0/6jlUixQ1i3Ykq50Q8jgmDH+PCgmoW48GKxugLW
SUamamXFI0WAcxMkDxxnTC65MtlDQM6IOPWpKAb7ZrjG2g8fUnbrEYe9+Axme8k3HWc5fh8pNtqn
mE6iU/evcLalZ+pALBXos246Ox7d/rxwPS+dGaxX4eySZmmoTx0gmeMmI0rvGSRwt3uugQXHWtaL
HElUSQoVK/H6fvuLe+2yhcAUUqfqcF8bBO5WJSEKefBsseyYwKxPipJMMpqHTtPmc29oFf85HEf0
2O8G6M5f6YP1FSjzTj48KPHrjXEdCbiJTOMM5bme+g92GOAoGipQgOfrd5Tu9LLdSMfsFlTe/g9p
XBMNsDOZlC7Si/eCDiDrl2/j5RCS/HZmrtymlKvy7ZtKnxUMzuuXYDiYPfzyzA2BlAC9YxTxuG5f
t1A5Kt/3HIYJk8U+ZW7k98ltPo9N0MVoJCwh74HNNPkDL9NOqrF73PqkIqw+X5HLRKJ2mpaJnj2W
yj8+Qnaq38eeV5K7qS//wLmctqPW0nFshnm3H+uetJ0KhBLPAxraYIIvCWibYkfkUixUrhsY/4Ub
duLaVrmzLoTGz6k7jrjwW1CAvJ38S+y1u9FIH80HuhaU3lwGyFlMvwGZ4OKayZ6jBQAt+0r9F4MH
rIVU9UQaaz0n3p0IyThGWP+NvJwMW0nX/LjR4ZDKigBhgZUTmvHDNkOxEbH9+8by+4Upca2tpd3A
KEHzRn+hSN+40do85M05ABBoHzIk+nqwgelPwt9afPs3WSdiilixfpDTiFWMpzww4EOvV8L9nDQP
210fR8nabApuM1XJM3ABDNgqeCN9Qnbz1Jx5hj2wUABWjOtTqIU8XPvuIgF6mqpsxCYFZ5GrLKfd
40vVOoKP/0eTgKhQGRc80THuefcWIleWbypc+xvaImeqzNVaMi6fd4nBsVXv8GLghiJJsp2/Sot7
ezYt+EuM1oqmSIqFr4JuODGoPvGCQRXJWmfDO5vR/E76DMBOO6QgO5wo2r7XtiNFscjNQUCNPeC5
VyCJjXFcZT68vxO9VRbfMxj9nK8KxkdUAUfMLILfHHzTx0UsjuA1ORie/1lxpF7g0lPUHZBGsmCq
PQdYiCcaZWtgmTSQ2wOrV1g9H+foZCSmobZlUYIXI/Cp1K74DUwovS+IcrUJZczwzM8sEz8vGp+i
QL/CYBTyuxnJYBGuR6rbyEI2YEin3RTdB2UTzmk7D6RoKCZ8rPDEVz+il3zSrh62Zrgl2RV38rwJ
KNc2k2GhzN+3KXS5QX/XlDerSRWOvIVMjlfrLWxsU0LTeJwr6sTG4BVbLXCViU0Qx2ZcmqGadwrT
3yHnQKzv7hynToOsJJ1WEWTS+XrJRqRa9IrjDjjJ/6Cu0g5cAKs+/Ol3WYy1nMsVqlZ6xtZWGQxw
uYPM+kULwTk66N22PACSXBfdcblACPVwZGA0Ap0ESXUgq6if5KMG6Mf1eiTIaP0DY7U9uYp0dnIy
+vo3jtJC883W80cfl+WGZiKZoTycljs0/a2Qdm3HoIQVQzpOjCHC52hAllkZhKvjQ52aZMOg5VyM
zVh67Kyp03YxcZdPW7OEmgSAZAwSY+di2gzY9Dlccywbh6r8DBNPocS0tV9yfTBg130PfS8DACaU
RU5ng5fPk0f+KzfP5M6eLc1zBi5PeKTYiVL8SMhkPmTnUGgmBCI7N+VtLa4QpCcvmC0AVg+dyb8V
Jae/t4UhHXYIA4zMUniL+7Osss5li67rSv27VlPcEyWlcTo/1DTXCpEfCw/52P4VEsjItHXbInwQ
VnuA/RK2Gy+YCrvfZG9Z2Q8re9qVA7Vs0mt4pmigd9GSIzJ5/2Nfo/pCp749nwUBA1UCO2KDwKBP
tfbRd8bxx3kjoaVedWPKjUd4QLBgZIj9YsdxAuNt+heWBjdGA3KOYoGUJ/1Oa6/x71hn8TB8ojey
2Ktkt06gKNdemwuZL0WSMDNuq1zWBexTApDIdgQpfK/qnyJJKnWocnVTdJ1OIQH7VKEMXhnv5Bii
6YLmJP9OrgrXbOqiuN+jX1avYTayW3rvOamUnwh2ifXJdmG4Ry1RPIOSURCOG/QfWv788ffvolGe
0vTz4xiWVgL/NAPbg6RPlffpyINCfqz1BDI8KS8rFTvlqJ8GhkRFKmt9efU7ChckV6nVHtBDT1uQ
wqCjBAxcEoaO1DHmmarAv0cM91T8LkKiA+IUIrziHyjeHoNwdrkLaRUrALOxWxRVXqwRnMwNzdzW
1GaUs9DWLjV3nuDM6rdVLWh5iAm6L6nPzEYCrGMnjZ7lophZDDn/Qs/AL4vxBlSyi2GN01ocPAQ/
NSpq0aCFkYGoOa+tkDA4cYevsXyii9WQyQdb5xlhly9thAf7XGX1cnFI7fm+vO50PdAJqYo7c469
UJVNOPZVqb1YHbOTxTdQwyh2yhpxJhpSkyls+56tqCAZaVJQunA/tN5A27B5IyVKaLsQKrOC7a9m
1xdTMxHPreznnFZMKDHUO5b+czs3obSLPNIergYSpPLmJLYE0g4OfhmDWixcUA8Kiqd9qe+i6if6
zUgGfOdzoEIMnoMUAr6yCXbWWN2lhWyqLPxTIY/PH+jtG40LUUdPbORakSS2Y/McR0U/aydLZf/3
TDZjawPfSIfEjcJdn4KZNlxFKXB++fiAO9M9Lmq4IaEMQIZ2wnGeNG8xFsklQvipeOAMWsQ7+XtE
nKk8x1VD7qbPUENhPTuyhhuvjCOxIgpdQLHPhs+Pn0V/uxG77EkPRHJHLjqkItemXhXpMwY39+or
0F0AktuxNHFxGU6nkw/K3PntDtG1PVG+1mnBQWjn4HbRS7m6utwvHN4oM2YM/UcFbzvtkrk9iNMh
acBQoGjAXSZOdX8xeJyFhG8H7RkNJUHYFifkstFjwS56G7OUHMilvMSM0ok+rdpQezCvPeZvbM+y
lKQVmuj1qX+eDjSuUtUJ73zUfGS1TWGA00iFxAwUJ/CqYyk/s1WbJlnvf9HtCEuNK0kT1/xckcQJ
DgAhXtaWA17dRGbpuQ/dh3TH5NaFrhjVxUzSYzp+IzLSvwxF48RnbB0jAL9G+zBAa5Kp4KNB6qOi
3+RXPAgxfcv8CXzOiOXkSF6/4Q7zQmxnLZ7Y7AzrhZQIRnxoSwiTrSUojqG2tktnHEsbU+GaZdqb
PpM7uScGpQbqd2QbVrmr+K3XDSGxI+8Ic7hVmtkwBljJFvFkDJrgFmuxug022ZrMeRvwg3RdRcyX
t8fRnpcB54v1M7uEJEREvAypDKKJRZ8TZ74/E85N2AnZmn7hmhWq0H7kpToTvvT3aJ7oRcaus1gj
obdOeOPLQTBIakhRz+E//ipU7N+mGRcKB54xLCKdN9GnKLC/kKipQiBChITo/MULH23cThFRaNvD
7Spt6vagAnkJHjmhLu+31jHfdPR3EKMapIuCbAo9Il8nrIDBfk61PfezpfUeE8Apvc5ZMYi9zxzo
tJaGAWpjnUXXyUqfcEceetQvC1uWiQpLpK//RB94Tv+5hd33aCc7Zh/9Efg0PU4IEdhTHAdLKilj
UmN/DaC7oJ94OumEqqkXV/LcvoNvNzUe8dlIigRzYP3UKnoYtpvMdmUUXmEyUStfaPX2/nXVEBBe
LhNGwh3Rfm7/xmZ9isCat3gUoMmuOMVC6NQSb/eiZj/uSCkcJHmYsYQZV+b6a3p8dSC/cRD2KVyq
EFLzItUO/UnMgScsQ95SG+l6dYZckzNSBzuzC4w+F8npV7BepGsG9gVff58ODjDtVSjWoit6mX76
4N2eyiv9F7EDFl8M5v6h/lkMnw4LG6HVVmbxTUxpAm/1NcTm9pPQhMVJtuEJYxCu35t7GUHRtnDY
aLs7Q45arnSzrlwKH+/EtUQcMDz9zpDoJN+Uo0W2/cIUuWoGEm9PqSFT4afY7eqz6FDv1o5E4qSN
2CmIf7gNrtlHI8tr53FZ+bGrS76CO/87VKdDo9Fm5naar5CWhIX2JkP5JlwdEKTPL8Z8poiLUU5R
AAS2AuEHWetkd8Rr1Qs5S6UJtwd2JVFis4rBMpvL8fYUyhCwMNteSFuSZXOzTk6/CQSUDCzhFioe
NkhAac0coiEARD0FteBRvWr26uqwZMVRTbj9zoIi8FD7YJhrpBAu/D1BWWuhGvtRqBbIDaZFs2gg
2/loych2aUTdcitdvXpWnsUE2UwuVR4VvnfF5c6iQIDjddsFFPw25qo39+jIGRJtVl3f5vM0e/IE
XZU4u5Abns5tbvpK5AmQKS0w2M2F3mgqIm1ARNU/c0E3zWgYKhwFMNWMme9LNSaRX3Q8IdjCFD/c
WO83YADJpyUaeuX7elE2bE9OTJakoBzm1C+ePAoIrEzUvn5nSX61AhszrxP1zxgtHj3PHJFgCsi8
xT8/HUervLeyGhZn6tdwM5lZY5A7xjqmjqBd5CGlWTe/OlJv/+dNqX0RWJ+kR7zH4RITAZEeM7w6
qOqldBWkqB4ZoCPrfOlV4TqT7GRTQ2DfVpoYodI67KLqFuER6CQlTVCpZju+75tAUWKqRyMkyz8Z
XNK0VOSj0tKxR+FyGpUupEqYUwlSXSjUxoQL1bUz8SYS35Hzz1zTa70y5M1nL1vf9kbWJYwmbl4I
mC84J/WxEI7dwRKPrfjGoZlZ00waOqqmUwQT3yWXX59B6162+I2hWimz6gmo4rHH4APtScC0eOZc
xqQpjmjca4w1ACjPLp9WXIyDLexYRFBIC5qfVSZHfoWMT9+Hm+Yykj+xA6B3sGL2/4pCoaImUiQ6
Rxn1CDzrQCDngNAspLtoWC3l1DJ76leVkmvy/vhRmnSylTRM7sfK3SOL8nD6rsV4YLbkFFO2eZKg
sE79r2Z6qeFGolOBtdABoB7902JGgC1xHCUg02XyanHqtHxGy9XTFAbNR2DmkbiXz6GPIvK2xslg
KP63zAHLZMt+ua+1nCNUELz9e/V7d4j0oUi2PzjryXxy4cm1/SpMycuwV+7CzctPsriKOgcyLxj4
Tevt7SUO74HyIRaKprkocQyGzOQ0lnrlYKlCr5YCQyB9sEPzaNXPGzvClZKkCMIibJhrb07goRbd
p2kZLHbHcgFTeH4aXbSOVW+7H5iDJhkt/eYn+fO3u5RO2nrcfT7Qv9CkpwFqHgU8+VB5ofq+L4C3
oSYVf5g65bKBVqbfGIMWezbI6yrWLDIi0Ch4VtusqT7iRXTVOzLkNeg3gNH5QjdPD/vkYATaFYk4
CPQdOQWSwfh3NHRA4lpEGFSBiUwi81V9p7ZqZ5pBeSMrMWsI4nSoq3WKSIeZRgPOKJ5BKdWgonY4
HtaaaLhqFNMD3rrl6GDY+IStG54SzOgvXg/1ctOnYAmxV23vZHCqxY4V7lrXJBBarv3nULUI0xbu
418mobKyn+3R2B1j0xMC5DkYsFeFHfbcguVPL+Txkf3pUG+T3C9fpiDjZL9deN87woxu1ql2Fhai
OsjlZ40pW8ys/LsVMJumDGuWpQvrFztpXJRAN2WjMV8+7iLo9sHDwLToidmQRxR5MCHyx52BtyGB
tAxtSETH9PHgImi/b2fBPrg9rCenq+7IE7C5OjUylGc5hA8KnylrUyALJYsENbC+NxRCUdO5IBl7
EbH2itjWRJP8cCpHuB4FJWG0OcyuC8zDuuvAdE6+QaVUyXrkvzbG208dzps8isLesI8YQZdx8N+q
GJ79bV0SOmkuIG6qUKtOiqDDucCuVDvX2AbbY8TiJR6sIdqUCYY70ZRRRgZtDYCdMKfpIA5RvZ29
G+sfDIMYCblBYRWnwjbUp6PLIrrbrDcIELFzFkYI4dCaYsQXohkZ1g4uNJXnjPZIuJmyXLkwvXhv
e7bw1BO0F4cdVQyGER7vI2CKIYr+ZHP1RYLxFbh5Ygpez6661NcAAnRS5UwF4+9Fao3hAir560T0
1p/Cnk5824dKHacbj1kXp+VlFzjd9XzsW7z4IsmUyOqx9ZF+wxGppm6R9BxaUM5KGD2aK6JVIWxJ
TcKNZdvptfOxRgJOwlpEJVqAsyABm9DMteVB3Q7FWPt+Pov6mehExV8MezkgWVaUGaBEm8K0zX2r
ZV4jvXcnGKhWz1ymIS92ABs/AwXneWNV2O02PjKDPP7wCnbvdbJjat7QoSaIhCVcZ5V1+86WIcS8
8BNcOceib1f5x0/Rt/Z3+8hYSRKHWZp1wEMOFPwGHuinzBQhTRmfmSjGhR4nvF1LFvYy53hKon1v
5PO1Pi6rLMdKZc6EPJHDPfEShKDE2tE4TiVGbVX2VwEPj0e+sy9JXBlzNodHxzU3CdzPPJkCyA7W
cIqH0gQ0llA98IiAf4VPtlgcEovb8GefyR2luET3rtGGctZNHlZGbtEeaADhIY/kftl4X2lCs+d5
pE2LXD7/RNvZ/T2+uNlYDtt/8wQp85joYlCaoAtiSNuhNdRl6M2pESFsCDp5vtrXxEOjN2xMN9jJ
xa7YokUBBlpuPQGeTsfzE5a9aDJ3RNaO84avhzvIeDh7rQk+/5QD+GdPrm3seVM6QESOGD/k5rae
7EhGlo0gSAy4sGXmo089nkNholV/D5df7gpSB1XdfhwIBZVDBtEzGV+8LpRPY5MGyubBc3e7TAdb
d4c97tik2qmFUbMKqzQ4aHZAwD/4a1LgvvQYorYxIzM1LgTIx9YmbTYlc4jrUEGRRcKzf4YzQduH
uNwL74hP1eLSrMgep2LZjRcNvPEEMxMKCjOYwQ85xi8fA/2RT+hgT2V066lPgE50ko9+NCB3T2qB
LmOAjWgkV1BFAaSKpnUVSLKMhbxE1E60tDulazsmAa95nVoykZcKhlwLJcqEj4qaRuXx+VKW9R4M
H/W/rKLnxJFTkMR1D93xBKHvkqSnOevhCkxM4HL466nw2thZ9bajYwpza/73U/d8KxKuXm6lZuLO
/Df4D37QS9N+fDwqSPVTIRll7MrPjzmsPYMbWBvZAnQJ3heud/MCPE5Ac4VsU+MLUSrsgFYW48HE
0lJARp9GOs/Ta+NhZJykGcWm7XqkbacTJO/lIu+x5L1a+pSOSA5bfvsdZZkKIbandF7+948hGvf+
UnnAmyVRWF8r5rVtiZG6VBSNbbU5g7WuI0BECD20xFJVMru4s+0y63vett7XpDcpxTQOp+OXQ5y9
hX5AqoYgBMgNtKy3FUzjn91BQ/qIfCYxqtLCo+uFh1JyceCQ7yD5odxwTHWL9BmO6KEj2Q8DnaSl
VBRJYomaqFQtnlcq/WOiKBj5b3e/7Q4l8wQCb/71isxzxa4rIGnvrtloeTGduUnMvcCIViajfJYE
6RyToy5XM0A6Y7DDLSROv5b0bCBh4jAtwbUUNM2j0M7yGlZ/NdpMRIiIqUptDEkOv55a5OuY5k+M
z5qKnGrbdieyorlPK3QjTWpSTbFgtxetpBGXPori9rP0f3CXh8Bk7aqicAVOlOWPi8H3D+bdSSFw
Q80dNwoOURwsc+PiN7td8nZr/qSzjto4GbMmSyiYXd3QkyOvwT1P+jywxFZJLl3NYoBLz114bMH7
fjJat/19vU8JQO0MAuBDKDrSQZQQjDx3xgINakcModNJFuHmUD9g3E46wAOSbOORn0efN0JRoV48
NrfEQcOGDgm1oj9+dTU1pi63xGov8iskRAMhqz30Z2K+6zMDc9TwIWN8JmqONh3xAqkfpnQX4Uqn
vk1t/uv412zBzAUnJrC7HMr7aB/My25DPdrjMWAMerXI2SpZ5FfFtK40G2lKbiNoTNm5PYiKHqm5
EyBEXCB0yeRRRkEXtD/WHFtqWEjWP78XcCbLHzGl4+rLPDcBNeISjsiDq6oWdZNmvkC2/iCvHeoX
OSBKcofO1hpnDdNbCMfeddi4xcxYGfFuSazq/8zbVDQJC7F4KilR6mkj0wSaJV69T6dUHV5X3ltk
Qs3a+wpt/jP6Ax2RWgYH3hiPY8/6ji3pTCsfb/40avAuRn0AY9p6jGR+SmDiHrwgEBY5j9CqImcf
EeiFjbIed9wZdYGN8SBbGNlJ9SlvqaQ/qapFSFBwAdMMj6KHhN0KAamlj4duO+tz4Bj5x76tRTcj
IHifvZDPT5PHHUvMP/1cN5xdh71d93xOkB93IQYuASfgPQsBQV4pP9y6Z74j6k6dlG17JGp8V+zv
sFKa5Or2Bv/Vsr2PNjedq4RqgBwC+YcSx6fw8W0TfA5qFySuVxLJJC3htYwRu4GhZUIx85JWorbH
zdU+1eRxX1/vCkpyMw45azykqPZx/47p380qrJfrhNLi84ypeH0MqM+QIqNq6uKdmhgqIZH0mAt1
sLf0xxFvCMKqyP9Eh3rrB+Xa/++8GtfFHggnafWr4mGzzEutrz1HjwntkQ4rpWbXPgULCEbs1wqj
tDAjQXJFpjHuGyxA3N8sAnmY1TbyxBCAE5l8m6l4+OgnVgEDE7+9V6s1/aTDFlThu+Kh8BWckNQI
ox4eS4SydSWLsRiQdqkZwX0sW82xtS7CIzecoolY5q3sFd0nUFMWar2rcsmEAWGU/ZaZiRP82c+5
OOW5CXY8AEYvlaWjomLiswDFwimpnTXq2Pbz0rDX7UKalqPly6OG83qxR/WFMOOk7nZji3MCiun5
Bsx3ADBDYLKhrBAT2JPUoSoutA45h4xQqV+H44EUOd1HO5Ok9y08SIR0kRMwRUa7EF9jTATEPtTm
kVjoJCiaNXI+VdN5vVbDtBZ4GDoQgCKuLUNAd9qdzLnzXWcxSR2+YYn7CnW0o7FhQVY3JNLyepnB
Sy1/cTcESUTjUY0JH4KsP0KybyoCGyRRT8Nyvx6Z84JJzcqlv/89ZyPGZctdkwVb60m9OQR1puiG
q33HrwtcOCYcm3eGommowYdeHybp6jgVA82HlF6cIHrxBKwYU7ZX5vk8KdUObaA38L1BQVWr31Vc
kttoDCaenc2r3kz25oiaWJYtKCZo2XgbMIvjOz6eLN1eEDtGeVpnwgkFLJ1peHO6fljeeJr+hPcj
gcAJJ2GgnTSvW2v4md3NTDpUYzGZior8pEo/Wzx+lqPND9A05Q3/zeYtx5VELYDDJ/4UYtj99LAb
MZiXU3qNKxs/qq6YMjU+FfV+ov5uaaACP+JZvKJy9Vy4zRZoAwdxvz/phlOmzmts6zCR28M078cX
SCkyZqE9ChD9CxbtgN4w0Ul+ttu+ct9A6h8UnDNbBpcvMqZqswRdyxSUC3N25D971fLOeXMACwxv
wfjLTw2/7niiMqQiwQg6aZDBvM8ORf1RciTxRj/wpxwh7WMMg5WeHbZ3zxn7iVStMbYquoK/BUk0
3RqcXhVF0sMYR04p/jVbFIvJPCn+InwxCXNLfTxbq40Y1modsdzoWco7tBvdYnCajv8m8ux9n7WO
vwF9uQiroLWWMppYGbLUHH8FDUQIA6WARSbJjUwaf352RbfvdEfS5vC2tXpQUOIY4kVlHNFS3rwU
VP4burkRX53fjEItXvfZaG5Nfu5OglNna+fvd3tJtuGoMLD6karSJtvJe+UAGpW+BRlVgNFr0xKv
PEqQJJQW4qMe0QRqG/gIbZhbjrPzyiAAdRbO4NsAmKdfDIbI1xD7Y67MWJWLb1yHbhV7VniK1OhT
aO+EhZToxISdlI/osw3gz3k38XCQYlpy9FEy7bH6BjVrBReZ0F5+QyarntMsi/rasqc6tbPNPuIw
EnsTkqNz2RR/mE3zaufG68AsXXDfmLhcJCPho9BlaFnvj9EGYlV2c+ieVdUwAjaS/PZ58dJFoJCj
LoVit06I4Ukw/OK8vMg194Gevd86MJkDROF4+AqGP8DHHCRl6bajWF5I9qHJjlBAckdEaYPPwyGp
PjCacz11sZybsTbTixNm4OLl/N+pZFCYfbhbjC7nZ3WVtZvpGDBua9qQPt2ZcGPbvKC12RzxpCFE
22tR3cSlhmJ+C6syj+1GMjBp9zx/3N5rQxsELUDp217KIqTYE8IxOVqjcO6TdrBcYd9aQtYiaEAo
f+V0vAdHGl20Emd3weDMbBDCp6mP+L34ZNqYKL1P06hoXRZxUgtfPZCILGY98q02jIrQ8DNXdVAR
ak3MXneowgRPFf7iJxwKoDKjzaF7JFAQNy6Qz/4jr0x6iNcG069V64QYGxSy3qoF+gsptjKFw9Zz
fcIaUlxZ45GZxR/k3KN9VuXCkeCZoqYvCz4wavdS6/CWZkpCuXMg1DJQQuWSnSV+aGoFZQQ9rr+p
1v9VuYhW97jYTJuSU8BAH71vdfjb2qUhH0Sb+zCbo2A+xEPmiX03k7CY0nacqDjZLRqVMn42/U2P
tQqWWESBRgUK1o5Qsa9kjyywx9Dydis1MNGVj3eHNirjpubgLocK8PP7qTO48us7P59qBHqpewUr
tTvrIhyZuP4LJkP0fEq/uW39Y2XBwDmshVLzqSitDWobet0gEcryxOGLr6dDlYtNysgiHtvPSMWK
ZSnrhfPU/MKLobJkbpjXmgN6eyYGOLrioAOlBiBjarNrlegL6hoBgaBbIH18f0NpqQIgpuUkn3gk
wzAZRJmyKMfW3e/rIKqCXKau+YfNmU+BPGItUw7ZykCpiZTkR+qc4MGpLlvOlHaFvzKTuKEqDMYX
T07LdgOAeQugngb/fgCvEwe4+1fzsajCimT0DrNfyzKmmFuf/Y/ES8MnNf3NXr14g8UJWZr6ID7p
jm+H+OqzdPzFjv6uJ4MB4wwbS2Ta0Nq4y01W60qNKnK715894wzOZJpwEH2alW/Cq54z3eKrJdB/
G/2fiD716eSCEkTvacgdV99vO4BzsuKwVLQz+TP1EdAhH1r5gKvwpKHBSnqJDyAdTsnnHt4c7G3J
Km5AomvSn/9Wg7+dQmcNs50Qr1AX8wFJdRcYzo6++Fiv9TJVYaN2qSSyTzzhuJJzP8rFApm744U3
IniCV20sQaAFRXN1pqwK+Wauu3O9rqUw3GfIFxYpaMdBDWgBMXMUoFCXmcAlLHW3k3yZGNbkOCNu
i4kpTdqQxK7+nJjeTtwMlDi0KIe7Sz1g1RjXiB7M/JwCFR63mmwG7FxDoJrCZV7xqVR2RVBh5k1S
xWMUGrVAb8GnkD5upJtRfbo98ahR6/dL2Fw5hp8rJZxGq0NjxEBB6nrCXlZUSYPjVPgKrVhQ1ifo
8A1nrKxTUfOvq5YjemZvOahWzOLAYfpei0XZNDpSuQQepYUceS7CGYwHpFKyDYjCUwElDhJiL+dj
sHZjH+XPX/7II6nBZBNy3r39sWPRBhNxweHE4OEnAoXjRfEOQ5uBDG/qLf23MAhpQ5+waFvDl+uB
1mN+0XV9yHUXVSa51jE04/IycGcOdtD/SWSF2nCsZLxGstnS+Tdcn08FLjros3lppd4mMW5oH5uS
ISsAuuErDdjAQxCoKSQswtK6V5imxmyG8MqLZMcPi6aMO5ZGnFiVMjEbO77x+zQ+4eDics0XZaCc
LsrnYRW4JfboTFdfXRAQEUNUMmVBSLx0v8+NgesjwebN3rakd+hh927r7sw6EwvfqVKi6UKw+8pQ
rDwrb9CtqMHqdjVk3yQvGyw/etb903hinPCDqzVaiLX0Vj4wzuDwnxC3Ck7SKZ6duppzWBlIaFdF
snkMsU8972uo7gfsKdOyzJa9qPMxiTBLzT5EbgD5lXtx2mPXyZRQIskVnbMegSGkLqKbiCPEZPIA
MZknS58RiKJrHPud5+qp011psqiA7B5ntdgMQQAr8w8AS2E3xtMQcAtlftA09Xoj9BGYAdsiHZsG
fe/pGoEI94OPh+qCZOZqtvQ3xZ83FXM+ve5vnoNYvY0j26/iCanLRF+Ntm0HOiQrEHQdMpQzJyJu
nuY2k6BleRGf194j9H4cOT5OX9iFC032w6KXEyGc9Xi3a/yuLaM1OBcuZDkPY5yZRcPfwPfIRLQ7
KBNYA2/lGzCPajAuntOAcQ5WYknKeYFCZuwPEX+hI6FhReGF01A48XQQ2CeAQTqa66c9h2smIpun
sCO9CRgGWwRGa4l3simK1EGXQ1wLj/OPDe48Wiix2pJunLlbT9/X/+fDqyp5cei3WlKAZCbUrxTm
hUiD56lsGpatAgG17fztDikhGZXg3dBaJCRWsMxCTHe4ik6+9R3ArI3CkLyWbxtwxXhvTHlUTh9d
4xvIJlA0rkpprP3jpFmlzGiMglh4ec9l2dq6c0wpwIw83k7DkoEXAgD5+WPvr9JNlilAlcxe0+UV
ydHTlrG2f6vAOQEWro5Ej97wroGZoDbz8AULeKxPmLVFzon8SIoz1okab1m/ZQghuI63BbfgXDqf
yvQRbcwPDZI487EqtW5MFqPG8JUDlF78YyPNx1mKvwcBvSaYlpIb505qs65XCJ7LqHLjtF2HReKn
85uUkxZ5jai3owVJdj75JwYpxCaCbfHpHecEE2xwr0jCnJjoDJGKSVzT5R1nLOrks+GmkJGysLEG
x/5JB/JHcTNnfGxhnHOKFv+cbtBI0qcYwN4gkxZ6zzBxnJ3tFksWVD9ZiITQP8+vby6aaJjt7oJG
lUECkngahiu8xJ6mS5hm0OnLmqk8iCfMIlDdWACGqBJURnECwQGXmU7m/AiqS+d9+Au+bis1pzgC
eD9YrfnK2xH+SDyhqYcM785tbMfq7PygNdYRa4J+55N0lPL8xVw6PhTwvtM5IGCIvGzCIT7ZbNfv
ptApt6kjdtIusEwhhpcid039c4U3N6QSkpD1ZPEvMkFxKhDNSoushhHqMsahBvLk++dIOGdoPChx
oUzDxKJctjdD13A5LCM7kZbDsdd4ivj5vLf9V1F3t6zNLtNdeYa1Q9GzMC/xV5DGK+5eJJoEoCLX
jNoeYZTlAlKUTpg35PeBMX4ykBjVlwkJOumCj2CpuL9bjLpXY2LHIBKFGaStkjU6JCcEjJqNChVo
swoGHDnP2OJDnEmbTVxgZr/ZwYKb+3A4Harg/bg1Z5BOrpXKkz+1f/TyFcKYGIU+hCln7b2pBS/G
seq5X1Ijcqqkig6/ca0kfW6nB+uVbydXLRe8o+tFRWJ/3zZC+hdwdec5QHowroucAauf6Mz6xGlq
twzTtbINPEbW5NTLhlNwUnRI/bi0y3lyY+59XSz6xAIiUkJG/baMmAIk3VCeJWanF0hUxsPiCfHf
hDipUS+bICMJ1HGEB4CTv7ekJY8qttYfOJmxcsAInzBJTllIMnhJUfblxTH6b74ssfH6TI7yjhqE
r6ePnFZSu8JT8m7CMTd+nZE0pGcdCR9qNLwhqVnjVTOGf14hnYFldHLkeq2BlYdZYfU7DL7UdEZt
MHYjZiMAuP6no3mssoQfQv8TcgYFjXwI1WACwtv19OzNj+AkpoT4IRAi6Ed6HJG7/pp+PSNZ9Car
j/RGFhUzUat6AiERiW5w7HEIm6jj1v6K9nwh24WF7GOe3CESK2lXiVyeLUSM5725fz/DPEmFoJBq
BT9aAAVB12NA1dMolVPP9rRWbUK38KwfW+DJKQGA5njgUy7zjpyYlmu9roW37UPxl1rzcxLSVdIM
rfPep+a7cW0pksIwym3MgEj1sLb+lpAMYDNz0deNgKsoxn2AnSDnyJJbkCzNFgxW1Z1Qhm7obSK8
vGkNtY4MesvVuyKBapI62KzPby1OFLrMVZ0TmFJNJetIV48dfdPCEtmJfZGQYWorzryFlmwdwEcO
YU3Jb2sLcEZMPR6PSe7H2sSq06KoW0RPnduiGS7KRkLEP6la7k5+FNu02ur24+y24YSygU934hoG
97oXOPwZ2Mt90z5yMQ6mV47Hhwp+WTGhi8HfcNhMknoSxtbw3pYHhCU0sBLXCfAPIGnIVuj4HxHU
OauSn40+Vj/ojpUbPjDiR/bpVbDqFe1tR99ruMYPJcm+y4JBXAKFNuq0uopRafIa6rHKqNpxOaKU
4zINmfyA9HTaGgThRrgGvN24VMCqBxJ3O1dWOw24LLi+A0TWLdSgI91Kc+h4I8yy4T91Xn1arrQe
/RZZbAVhDg0Gm+tuMKzFXPTN6EzoHAlYfADCPWUOkEkfrWgw0g+CqeJ5jFCui0gqm5wCbUAwVuI7
A+GGd9R6jcf+LYvZIRLbgiDuucIEhbF0DENXsbbemUPYtaNYj4lQcNSjLAy3qZKP+jrYD5bSPy0R
Eg7p4hMA5IbxrlsMxB6cmIpehkL1m9q83plOb8pMS/hjoR9wFH2uCINgNSPjE2DNp8A1M4nHWFXE
O5OR8O5nK0f9Ufna+cI7npibO1NUzPZMmMAwwMdQ6Lh2xlQJUmXz50EQhc2QMgAhHWC7GQIR1mf2
WZEyDUmGhoc5KtayIvTjBSDe4/GsFOWJaAHiTs3+YqbVhyaNKCiVKvOak75gW89pfpls+A/X4UcR
ydoFWz5+7unHHaiKkXdiYe6W/YqY8JYYn4W58urIRa4HWNtFsAnNtg9mWWyu7MYQkwfUH+jZx+ED
Kd+QCiuZy09yqInkarvzpS12DsyOVvTFWENdfNiXlEvWnY0qUguykzr6wakprFptboBv5kRRFwU0
nkgNqgvf7EJNCMbKEjr7Gooqh1BJgLwg95HDfmggYpJVAww0zuW6pMdTkkX1Cc5+jr9Q3H/9EJYE
uLEWqCtp2YyViENCt8jDNd7HKjeC06rZsSCviV2dOc9MK7sAeQB/yGoAAHAER3jwbBEAg+00Hu4T
gd7FYsVoDJYLtPj8jHp1MU5Fk8hOxy3sUttkb49nnc7xU6jHjzJJYRVLcdbpF96Kc+4zgccMrdYr
J9oQl13zI8rtx9v0GwWIUnkQxE//d5UxjLHBpn6tDJrfkx8GsgpM9Up5AzHGStTYweKZFRrPXJu0
DHU6E8ZXQGn465wXpLgLDlphT/mZ+yRlBNzDHIbD6kSwgWWqeWbuZCpEozRNIu6zsh/CCyrxqQY8
7hyy8TnHl//Gz1SvR1VRP/M8xMH0DWsaXSItGgDrWeHEevcu+V4apVIk+X19Bim4T+nlQkCkqRg1
L8h3fDwwxCgS/aD4mCEDd4KScIzqb4u1aEtmgWgE2QUWlOOHyrBU/XRpcYiNPYHlOdriuZ7jULMN
J9FeGKng+59OqNUBiPY2Qcy+OSjz3MtkHkhm0O9Fh/gvz9uU5NUqZ1LKnZCFe3gFC4kQJ+zZMeAz
v4lCl5+ci7j9VtYrnhc5MuoDWVtw+YGP4Wp5yAxL3LhJ/LzrK8A2xAIHd/oEu+ki4+TrQ6wmh8og
u/lXEfRSkybuEE5B02bEQGkVmNyF6XAyy+2Wz42UehL41EXPOzlXQaNWGehRQS9UztPSO2eGQp+W
cuLVQy1LGJme47pcBiYiq3hTjW7HlyvJ5CLqf7++7gVwK7T5cSHAAVxCF2s59Kfl3qD676tpE5Cw
Te79COqQ2td2rGGNWEFAji10pJqVm5OxhenRRlXfAtBzXOiNzv+RAVUB7HfDaU47G7LcuOtLp+RV
tGb/xvkkgg41CGMKyninxfI6UNjHROvSEgRYn87evF7+lyiZ+lKglU1aW19l3KDP6aAprmQ9Kka4
3suoqwYL6Bkrea+FMKhKbtdhtFTtf2aS/NcyAVctHN86w2Fzh51ajSaCZfiB7ChVlvgTU55wkduj
ljdRBiqrEcaZwMlJhW2W3ExEpJdxI8smAlQmwYjQzcd8JDvEwHRtsAT7aHZWTzRxLAUhu7KlpotU
buK43rGa/NLMJwLErYoxPIiWOBzqKDxbkMCs8xltsh3O26BBKM0bNmejf3JU0vFaxRXXwX5MPAt1
WMpAWocVqkXVVKuEjuGdT/WcCc3Zj6+ozivLQiiv0b2gZmG5mWGIqaByB2ydKV2G8vhsbQXewznW
EqZwMp8q0ErkN8vGbmF6JFtfeWnhgVels9no2g98YKM1kd2bXJkDgfV35cOVS6/w2ejdKei7Ub9J
9J0Y0x/e+PSENgBCi6LSwyjcN5iXSEk1O3jF7igAno2HDUDBKEQJ6qulnXl48y8x/GwgbAKfvCpX
b2oCCRRutOKpm0D0Bvwy6rr6apmvDSd+2aiwjdaOV8Pl4ObGW60H3i83t/q9KvPCzSsUplvZIcxW
uXXDdiDhFXL85L2qVaFoEw460C7mpWIKrA0XYa/3aYjHTtij1sFPVZNOKbKOFPZ/uYXyenqPL5fl
yYDMu5mDq2MAWOJmllwlmNkdCf7PQQKY/inZCxJjvg7ZmmkC8y6+vBvzhiATXeV236P6ALlGBRdB
UI9RAhSfq9cWDHNgGtmI/NieDOkC7bxmN0TjyMuZ8c5Tl4WUa8buo+D4cUT8JDGDc0rxTxTb0Evi
KVl+RLu6xis10/FRwgkAWJ8zRecSWwWqBPnFwl8avJZGdp394xaLXTxVRiPf7pPR/zreQGcQt4L5
kDLkgMM/EuaZaa1D1v5cZi09a2+oDXiH6u6q/LV46cdMykch3I3wfTj5qQJx8inFFlIDl97CONKt
1YItUFEFfPZMHHY076EAlwBquXrFUPhlucXeGs78yTIxPAN75wllfYjNuzM4tPml+VxXl5A0RET2
+W18JvgUyB4OFiwKjqexUTPbDNsaadPEPdU5UyV14kKH21FKc4zOcwcil88RGatX04q5kffnOXNj
O8xRMghTT+1vwMP/+tuuCCftxDFVw+NnqUQkafNfmv4EWgEl0pyCwZV2eprTn3+P2NUnbH6BmmFn
Zia4l7idwGHOKiCyqrV7VOhFR8zmksX0YlweEAe9cWm0JyFsRsNJ/3NWTIxOJqEWOhKoy/RZaGrC
8SgcjdaQ0zztIAkjNoCuYWeXGj4oBPQnENHy8GeQYgGOG0omX4Ruw/AozXMV2cN51CJJQO7fJOT4
ZkLs5BGCCmC8auTvM/7h+AubP5UtRUjrF+eMR5LOoP+6yFcO09rZteGqGrN0Ab7/g7tq4+jMsDJZ
sBllE23VAxpN+EhOdQ+8Dp+ACV3KAHE0hf/9RZRhvwZ73wpdC/kmu2uQZMLkT1qhwhNMvJWvoA6J
J0kgsLLL421dk5vXTsznTsfTJbqh8QorzXbjtltLbH22403DbFyqeQdDpcQZMvdc7wftDuDiwAZr
HGIMidLf/UiOzZur4Hl+9q4dvcLezojunQk0BlNeDWuFKk0DfSGPCfG9iUnvEjxCbBzJmNcSF7vU
n7La/lcu7ZtKaBfGIw0yUP49fLUFCHxdNOohlPxxTToVFisPhydpNTmVXVjL84UpPTMc04URgqU2
u4Smwq2CmvLU21tTui+HAfky0W6zd+c8Q2Qhqpzqcg8/bPNvaxI9TSR2N0LAN5+hrGoPP8ESTNPi
FR70XGEDhuf6QMl8W/xLZzUR+9KoUKFmLwpJWJwVnHEJ10vO8CluaUPSlI/2VoUEjC45TVxGjj5o
ZMS8qPMB/1epivnxd0FL2dEZVwVPFokcjHCcToSFO6X/jfltgijYRLyOPqLio+5g9RpnMVFXkPg9
JOaxhvxmM6ac87Y2a0rqpwS9qLS6Y89ZkPQL5g5ndNXsm0UJ9JzReFe90BJg2G6DXZW0L67+2+Hj
q9aQ79Bcl5h4zSlwZUHSlgdQSDUvI0CLWU1Z9ireqcuKASozl44sDPayZfr/yJI2ZE3cdIbdsl5O
1Ep1UTiN7xjcbI6Gvn9OhdhDJJm/htvJp0/emjwMAAXTlUFlWZ4s42i+SHzTvNuekbnwdGbXX+KY
0rGMtaN24IDhAvenKYz2M+ZcjNAq4inQTDDuOwGZLskmNQKIban3vduUNI/9KMWJZnbQrccVK+M6
egIisAU6I1otTLwA3xf6nuqKe9qyK8c1hvscIB0HFQWByxgQPrUcV5Uyn4ZI1Vhifg+uPh79B1Du
K7kAe9d5aeDyNAEsWMhuEd/dCtK2HPq/Ipsv7YsghODkSkuSxofFM8SjhoEKMMoP13rT8haaeVh9
llYUYO9QXsQmIAtxOc+w0EjNDJbKxMWDZnILh2J0UEn3DOm+U/ShnST6XyemMk00b7HGozlsFVRk
UWLx7HXA13SVFF6k1AdFhq3Q+9KxV/q1+v1h15bR5NqD+TazO3UwkCks2Xk77OLWJHrPxvjhco2d
GzIKgp0aflVPYGNd7CUo7A56MVYTn2q6o6+iKupPc7Wo4p/yYWXtDlCE5dGkIVuQfM7PGEaao5Fx
T/BpwEfGQsdJL6Fs0fhPdyiqtrMG3Y4ft6cne2MhMFrdjNcM62s7K3MSD0r/R+uuPm7RDxK3ngiE
SFuBrVDJb+VqHg+6GgkA1IqSSOzs0EDcITls9iN/b9qV5dcYjb5XclxzNu8XfEW8dPDAJQzinSuF
5i2yIDc7caIPBJRfmCIHA01xFoRup4ccx8C9nrh+EThnx2f73ZZJXsy3+gt3OMiGTMV2phwRMb9q
a0ddxcpCoMemXOjv9Ch20S5nfgUAgecBCXzeho8wpotlgJd06JQSNsSm9XpEc5CLU/zdUpgY2sGH
sZfErgbcRRiHCE6KSF4onEguD41ois1xPkzd/QhnulwCwkRvcgbmPcvjGTi7v65qRAWcy/BJ319M
nOzQMVIAi4vT2mFhB2uK3x7GnaSTnHi54ZKUwLluU+STuoMAZNphtwG7pRxHdtRK/y6hdC9zSii4
flzcigc6uTrEOeWgT92fb4QmthF0MDzm5zLg+FcVdBhfRoXmrlw/9BLTuZn+NlMxupAYaHc75utt
h54jEQuRWNtiXiUOVSa9hCny9V7aJV/oSb8jeHjtaKV+wQjCEBCJJcW1h4utr8Ermt1uAvTkBvKC
gHmH+ZIfk2UhVccehYSxfnFagC1u7+eYnoVDuQ4tf+KfLI2LD1Ev1FjpUHNGOZy4bibRqGSKpa8f
D7busrkK986StxsbL2u+SAb4XILIU6h2vXG6KdeyiJ8uZEvIS6VoBgboqvbHIHBbxZUHml+8z23z
gxGByI3L8it//7CLMvVMAFLBEvgZa/uXQOnYiI2X1ZnR2/73rn4d37B3b02i7db7PKp2OcC4qfSe
vL3F53SC2IR37dzhYcgUv1S6TaZ4x67mOpAkG6QRHYPxskIfPTiTLgZkvGq6KQcenKcksqsWTVJC
Rx7H0waJgYm6OwaA5x2kPN8nqI0OhPCDtnAjSiAyUSFlzEZKhSC1UgrRCNqJ84LB1kg1914SaTun
dVbnVgr7U7AzZSmpaqChMCG2mPZHtyyxDGsY9qvx/UbTrw1G+OOJzDi24DS3lruFLMP0kcXbuxBs
PnxSmnKShDFtOj4SXR8zjq8PcsVaD9txiSExcS7hovm8xuFUZsIa7K/lBfmevWFpL47eL1qSooco
GoXm6WmjmarzP0eZpS2nWZjR75ZemwDSA54FRrtfAJVcqnezF4roDU5ZEkpn+rJ432t1Byd2roJa
A4xNWmknN1GUSI3edUf/FbI4fFK4U10X8W5PV6wVbFlzvMtG4ut5oSP73TvbrF7msrf5pUOVAxUW
0xbzJjA++AvZ8GEexcuIB+28dQ6aBdoO7R6jQeW+Z52yT2LCGby3bxIt+5BjDGdRB3r19q5IX8XW
Y4vGifDFq8etXRCxj2Mofomlkc7vR7L93CLn28ATKrGGF7tyRZ9rKQktMmiudcD9pLqoQoLhMHfo
iU+8Exnp6KMPVcATm1H7ob368d0S6DpjZuCTczZms8yubAoEB0FU18DfL+nxHHBv5m2CCpIRlKmF
hPV0x7IXxr/xWJU2fcY9gZZfkasQDB9mFWxhH5xFaijgIwSv2NNhvAT1g8po7NXXPLIc0M/uUZsP
rtnyLIfrwP3n4g8tu5xhFPud+yuBzEhEqvAefohXYfcm76b/VvF5titQ0YUWB7I7tzxExCTutJoP
Rci23GeeL4CdXokZ4eaYGjzoFopM7KPcoUMgKXgF8TYPd6vdQSqgVf5/4sUsTD792OILOsGrla3A
uAtEcNeMu7gOnq08xNNARMYx4W5VSUfSq6lQXFjuma8+GhYl+WINSV+s9ShLe04OXb5+MZZqkB8X
lwh6lAUefWOxojxDQyEiV+kxSN6UyT44TcCA0NARKRPguch0Nf9uLVqOObDIpxXhKjJhLwkST8UI
YEhnj+/j9ntFrA+ETT/MtXxsmCKJj6EvbATyBhinA9pn+rL3BGoUXo2/550afakHBM6CvbvcxzHf
7beSCfxu5OTJgXvfRqb0+LtOVd95NArr0KOuw6VP5+nSm7R9sMy5Hod9+N2o0aOCmcArBI8frMQY
+ddeHyZ8vvMbkDuTo8RTNH6ZakR3nw3Jj8+AHSFBAnyv/7jAwPi8aQ6lQ90fsXL/oyLau8z2cnlV
twNn4KJqSc7TfZXuivGCa6bGYXa1aJwqocbPzG3BY5H/EusNOi8ix41aoQ40BbyEJ9iBjgJyarKj
OsOKt8xaDC7XCEKZSsyHNQqrgKlJwm9h3f4dszR8kLNZsDgr3YVeUrK8zZHNjsDg33wE1qBcZEBv
vUfTYpGI5vJIrKd4xu+aypsdnJ+quhyVm96DNrOY4hHqBpS3Lt8DCJNT11CylEiJ7+KqQD3veqoM
5L6gB1T1qx3NGw0KqJoseFw8YhG7DeV09V5E0rrru1xh7/MMngV8d2TgiVqaSPqEr44GvXrZTwME
e4PNU5fIDlqtEGQ6gBPmYzoP1y2mxvOB3Zb5lWThRzhqcUKO/AcWcvnR22O9jDouUi9NiZejzhoU
095qEp5725rfY/8g2lVA0ZTlJFPW3l32IP8MuMZUtJD8tGpEMwiE0xxGtKfgGGZ1wkmSI+5fLT2I
kF5ndS82AirzVK/RtccHoRKN+x3huxTdOu3h1CWN6COL7ZnYDjePhgad2e7K4J1bxDfhX8heCMGG
Wea7lm6/pLB6h6D7tcQ4P6DDek7DnjPnVFNylruJVM/tAD3SbI7+rY/6LqNIFbjsNvF5ZFVBM7oI
JM7wB8fRzPB1ZsiMSfSKmcv1M5VsVrnsxj2ePa9uNZzvhc3bBoDxp8CBEmT/s4sAniOiLksf/A64
0NH8OpYD23yfXej0Ko8AlHtspNCTwncP5rwmw5p1LMG3TLBMpAvbNU4r4cbWn/tS2RdGSMmREXIu
ecqZtgGUQNZ9WB72VeB1KJfavs9rmkOqcu5uxKLiGeuCH49h3V+wqShDqbMGgz2yfxJ7m4sDEGzs
RZob3LUUh8lDXHI4ZX7radkAih26v+wneATxJuhqqQcRioN961ULUb+EqITLEUm7ONIMUilvtE2a
ykzL5dagRLkOQLNbZyrifdShSjPLP2XwI8EBw0eiBI084M/uX5HZCEEEZTAN7ZJ+eT+pgq1OD+z/
aRPnQs3RHO/LupzECxMzkjLzjFz2G17+UxWlFOoWTBwCCresosTbgP+Ga/TZTHqGfJPjiE+xr0pb
IVt4wRlrp7YuRd7YuntNUn560z4Pk8Mjy/KVjiWv7xnx04T9IWN9l7h9Utj6rof6t5dyHC/ubpTy
C8OTvmrrW0zabT6ih6iS+IG/kO0pWW3imxFprpoamjeP+irFc9OQ7zpYtOeZyl6LhDT1oPEwQYB+
ljsqSFm609WILIkpJE+aHXJwE+euM+oOFvlF9Wdq++ATpIo/gHcfciJAoDDPwqqGwv8DRuSkohxR
2CBSsY6fxJCWSz7+BVSCpgrFV5ZHIoMm+TA++Bh/BmQVFGRKKKLtouEX3ZEfHHfq8kE1sW6Q+KLB
brKzfdmDnfCcLVHmPtE8cM1KX45nsNvGKC//9OFzL9uXyjO3+gfbKwFirh5WWf/0NNcv6DXXfwj0
WJYAP1yHUsUJG9B4C7eltnHek89wcWxaRW8etzB10ZG9x9nRIMZa8inj+Vl12K7aAA6UnKLr39cK
eBtlfkKzcQNb93wWermNAMdiRDNUp6Hvgbzg5Shp/hmPqaCcsydS7eSujXA7wk/4MkNn+X7ZC0Bq
NZDw8tL/IxD2fDHQSE6l1LAge88XSVMct5rE/IAnKpPINNdR6cb2qqzZtyVK0r5J4w/6alcylpSe
qm0ffmf3R+DnviaoiXMs+WL7K4h1j0UWCdJFgq6ZagQwWUUIDvhdoBfFPzR2a31fbt5k+7GgT7xe
D4vzA91/xgvmlfY6HKBSHnFDAG4TbQ+q4sFEVak8oCXEfVnPrZPQ31VXzfrPNpAuzveyA8MX8d33
yuH07UhwfborXt6NEOvF0TXo90lP7XD1fawEYTbp3Ip/lWpd/mb0JMSflDCUuPUAlX6jiCV0GkAo
N+kAB10YTO96i5K7pCwXvj5Cb36tVD50i1fnp5BcX0l7YV2x01loHPjpXSmS9dQGfjPsa4HnKNAM
xm14fSKUtAw7PD93MsWPKolLvBEK0fM8o6mOsyqKqNJ+efLe9SlnHYsUtTSZb30j0b56fZIkODQT
n5baPsNSi2bc4AwlTKzQX/L6UJFB3qW93JG189sTH9N3W+Whd1UJCiaepg+N2Ak7MBuYMIwdZ0SK
rANgAK81zdnLZI/IHp57dM4mehYtdfJE+QqpjPG1tafHqBIa2RtW9mXxajVM80Wn0Qvf1+CMWCjn
tyyDH6aCqL3RA+uyjy5+68VbaukchjNq9h9Nhb7bklh0EbLmiK3jbyaFr81PzBA1tlG3JfyJ4Izz
YlQCIMCiH1gry6urMedd8EWvIcpnWm+MmsWLHQBebB+MizoJE50N2xHow1kb564f6jNrZLJXCMs+
spwkL8b3LT+w8rDxQsH6tPV6+l1jRxDsdtrBBfy8hMuQXjIcLlRADkU/gLiock+flL9RUpTZl1nN
thJ0RJ56Qj6i4dwZRdDpRXF3r7ML0hKKCkueBrk7BT/QMGc0zVUFOHnTCJ2a+d4uabUG7JANsBTq
vWHHnMbCS/xPHwdLoDlI4je0WSz/zO+RvSMRYIAvEFcp3x+a8bB0OoUbdfy3Gxkou2Rxi90kfbj3
zGfLWdc+1tf+tngmsxgltZfnkiQVl2PBlVrOWfejli9vYmppHD0vLgg9V5hzXGVTK2zYPAgTIs74
Bn7QC/ZTSehmdM/sM7YarnUBGKyYpmK5CcE9FHnM1+E3sDCN0hmb+3vP8uyDgmdRN+XM/7sOtpFm
k3yVhL2uvunENRARBfo3hJsXZQzTnJkXIYno40Z/qV7Fh6ZYvvHXX2UTo4hSvwyqjAdztJ0qY/UY
SC3GObHo8dXUCc5/c33q1Q/vnLqmlm/hc+A42c/LQrdE1nRC23q/khs8U3ztZB4EaqhVjO3Fl1Rv
PCBWMzf4xcFWR136NO1PADUwwSGW57bfWZs47sCcmR8AOlHw/Yw3ENpdx8dxpn0VWfeZaEiu+Rb/
QNUgACWG1FGY0kC3LLJLcM+M6BncmkRN6w/b8tegIGFcSZNnJ/HOwPJY8dfeqiY5Cw0zy0rh2pJ+
k0gwe++n/fcVe03dLL9qF0oRSOh8FaksufRSExGJl/iCFxMNN5q5EOkEsfiNQxEA5p5Raa44tluy
Oluv1rLy5uSA/8/mS+ycJzeW3IrcVdHmyFnMdSpVkcNdgeXKRMK8puwe1/fWaKduWujmc9LkOClk
AGDSSB6br6o7x4cQ5/L+YHbhh6Yg9uKWTlrvWTCtPtm7xefFw0Iu3iSQfZ9+EmGQJ3Gin6Mu2DoE
Pn5Ub1UQbt01HDbk0yMGSC19x1epPxnkVOqTjYOJAdct38QS0n2tCtEoEOjZG73+icfBOwlTq7P9
Gx/7yAEi8cAAy67fU8K7EDHVUEDPH+0D4JlQsr9x+twhTLkt3hd4BCxAnGEd6a6+d4kRp2oQnovS
iMZ+qyjbMdQBiEh7T4mlYgq8d9aIib42itNfb0n+drilFVnYg36m8GzS6bCooFCibkzzTrqQveFf
UBvRjaIQBYgvbg14gZLtbQWKblEh+Jgno6XEYGoKXMj8IA7+jawn6692zMZwO4oqDBNSrvWhGT6w
XjtxFw6C1dlA53P9IF55UMyHBIayBV0d8zg9vRY/l8q52f0PWRyB+3hjU/sA9fCrsOgQSs9GMmWT
akerAzNcTlNaXDQSO5/omwsouw7LYN7GnV4jesJ4Z73PlhyI9SLyoaTvGwPUHfu4TleaWmP1Kv3P
yMpmgI1rWmiCZ/qi7Szvey7Dt+ipH2EyFXTQCYh/jSZpEMlpZdpr3eC/tvGtUgfTqdJWXbYm/hP4
1tXgasc4sA1o6nWxsH87AKocN6S454ed+EBmNdkD+hkDnBPx5KzyQOfAx+zoeqA9GNTHwFO9qdpq
WIH0x/aYzxuBJb/gWPGLjCe5krCf8LZLUSboVABln8tMm1TEy3grqNPLQslGSHw3yM3gHFJQtGWf
KwMMC22BIAeByxAkdlfRrHCD5UFCSyxGLQt6rwC016GFkVVFPvhX0u8YiIB1K/C5lHw+Sgo8MSbc
Ds8U4JouTkNyugBLGzREzxLC8cvg31ZLJA/X/fDeN3NZm1Y9iIN1uxxvMzEc3zO6Q524FW+rfy5L
7xxxC0HOLBLfZorS0Qe6Nz9JITtxj/pcl9sxCEEpcmWRLnH1891CPcRY6IoRz6T+xr5pCSPy5GDW
zi2elLU9AK0apIlOg2EkvGz+81Tu3S+7MKusTMay5LofY7pg18u5AA9dvoGJ0Ux+yLddKomPqfgu
LFg3CzN47XKQ1ReuwLrzl22ugnK/uwoCN+DGmcZjqjr8V4q8ms92OHsWsMjRox1ruYcZhgaZQsBo
qPjQzjSk/kh7WIJWj3zwgOacoNcXRpt9wF2PV72ULJEOqCgV+yEzC8utE/zXKxcgglVolhoeduyC
OA7ktc2r2XTHaJa6VNp8ZdtVpR4ehkmTvyu3SeieJfvJ0Ysx8Rn1YZarfDyXtIRkK9/nXJqc5IJy
7xLmaXeH9MWTmGodTTjRm6+CrwAyx/XvnF/OPN9+Q3Yu7X4v34dvmc6KjadEO4Hk/D0qxyZcIjfh
gq8+tZy/wS6De/ysNgL3Ai7x8KkY3oc6EV2GkFk7BZfCFWhAxLRT2wbQXLvkg6WTrpvkjLkCxMR9
zrHiddd58MMif2DbhHcC8w4ljV4i6DbFcrN8uzDFMu4vNv4hFMwmj35Ho2tAv7UHu9rU/SVjx1H/
wBHh0LD8GjPJ4kBnoz4b/2rplUQ/0rS3taV4XQOLr2v6fzLM74b/LlPZKCxywhKAz1nJOPHdmFFF
DKZdf3IzYS+2ohcdhTFLCzq1fuGAWp9r4ewe/GXqgtvx4hBZXJEJSF7OHW4E49NVC0PrK4Ms4tFV
Ql3rddLeWMGHXFVhNOH0grjvI5VTiJhPhVWfZ3tUCeDYI4aLhL6/8102ZxC42buouViIz4gkvuCy
E/8c+KzKj5dh7bMisst8FUyW/e/D86ezlRwA12nuHkqlpGfJT+VfNTW5oD2jcUDfrR8MTOaDh8fp
K6xYnIfJp6rXbXBWs9kDjfbwz30pfHQU4m2lTKWWAqeMYEneRl5cwHPOL22E9cT7BGqY1abEBE7d
UQCK3Ar6vvK6rh2rDIpBc3ynMTPcGhWjH3GcFs9cI63v3cEIj/KJSKOqIH3WeFfGtCRM5gX9+o8j
1YKQS4Rz/KAxiKfbo8QM/8mpDup7i1W0A3bycJYCniY3HV+tAdz99oavpZsZ9HOpfiD1CJBNqhlX
dNI0xyx6F3Dj5xUARm3csdtQ/9obTrACs1CDoYO4M6feCrwz8OMEaRjSnQYaXy/BYqUZ4Z/VKRTI
Z0CBopjJq08N9Hux4GKnQhAKUvDUoWxBkTL+mKWS7rLVCyL/PjVP1fINSnWT8tG2oFIW41wiw+T/
Q5RftdQRLAEpNAozJ8jQPoyvC8sVC65XN0sX6FwnLCB1sSh+4AujMdg5YUFCCqm/EQ7K0L915tSf
a2yA4LGgoKlWrsAEByYnjQvVZ/6gQrf2wV5tZr809SdnAY2UZFRouU7l0O/QzHTWMrU9M80eHRyv
heuvwcXj5UjXvsSDUtdluo9k3QAtbn8wEx6WiPZ1NNupu1VQpOWbQPHK9+9aXwVffgPW+eqWBfkN
qmwyWv2GM4gag53vzDkqatl6ImveKhnAzIjRY+9NcI9XIC0lC+PWwK1Ub17DosTvK5Y8g0cuekBd
SmphP12waP+EZnjxXZv2UeVoV5jWs4vciZtqfm6AP95tlP1YbmMBfrHgfZod/PHc5oAK3smT7awv
08tuoepS5xbEgB0xqNJPUSYHWMFr1FVWg9v7EmJjASNqQm5k3xkqAI5X1qBfkW2z/prZEc6kGtol
m9aPcqDs8MWLdd+HQKF0tX1ImRgnykm/n53PVDx1LDV6dfmLjiFU+dYi579mORHR6p5WHCm08Fq/
oFmIXQMSBB43o+1tON2fp3FwGQeGVT3aSpfX3zbpszNFMiN39zbXyqSO1TceJBJC9qAjrnuBbyLi
kGjooOEg17IlNVJMoMhP8kTvDZPwBXifkS7q5t/Bd+XWQqU0T/pNd5m9hPMyG0GThir+JGynuOvG
9E9womQwlIdQF2zEHbJ4oM1o4zMPC7nn/UDCO7FgUd92TI2TNSd3cLlhRMpuKpEF8HgUdPZg1679
E1cqZrBvURpYdJYqwTxakJXhNdkKegmloXsByusCr57i0urGNnSG1DzbjnO7qvN+JOioPGkT1aJa
pPfNM6FaB0K19YNxDHccM7m7v58C85hLjx+Q2fD/AJ2+zAeZOXFr88Y8NtS1IFun9YrukcWKEMFd
YGty7+EoMS+5rTp4LP5TH9jX6J56PGnbhtEGkkEhWx2t72RKuSHr0mB4EwVQa9fbKNKC06xBRxGi
2l1iP8CG17pHgV57/baXzPLtLKiw5BbclqjSP6xJG+xagNw/ixoNMZfY1/bbKuaczKhUuyUSeuAY
BwA31iOlU5gIaiIr74tw+sfoDRePsthmiIEbLI3ZXwwZqVCDfWXNVlxrwAZNrkvF6RSz2dxOPQ5j
qzkUjBuiG+FmpgY3q4EGNiYP+73dHLA95+mdSk9/+8gvDQwYvrGAeGvXvX43B5IFI0rVgQkdtijY
PSPyBonGjj4FCj9csLEtvLiomIwjwI8QCQ9+fNJmQZj727iLMNmNGAV2r6iIx1dDQxQXVxWRen8D
hOvBWLchZdLz4jyGDK1aPoGBc9bjrK8e9Xn1j11ZWmLkCfbvDBhBzqRw9zMzmBmzoXWLhUrNh6cN
xYnBsDPnd1LKtjdPEPWRjtPQGhklxxkN5cn5vf72XxHtcXDj8INCErAwKXreZ7vdRmxPOj5cC3nh
T7rmTXN1T3QEQRY4adNk4ZgyujcA4R9SS2j9mrIGYhMgoVw402e8oyxbAqDXmnWe2YSMoYnQTqfT
GbrX/cp1EbxyDGSEsN0wOuDoq2xmotKoG22KqYoDF8ANpuAOGlK/9YdJv3fdRD21EZs9gr3Riaem
ZtqLxhNnuXjBU8YxkKWck5dz77h0ggCzULsCF8RLzz7GYIxg1YArCtmcdFuuWi92c6MuvK+f5fnQ
cnEx0VZ+Eb00smfZ4GPMfuWQDQ7j72z8QBTAq48GdPPbJBW5id0uIytXJkTFA9lC846kzPIeqC08
C57ssjEiriKT54eM34fHN2pOYGDMoF1hXtMIRdiqSkmCcsitF93IYDmtVjRPXbNrCvEtl847c6I6
gDLtvwBHizS4JXeV6k8NpYoLjx8CINH/hKCz+vVWWPyoeTuQBnFbtbEKwIMmyOCe03lvpIgD9BnJ
lj/ix/6qmqOpTtqQAOs8Qt4QSo4QwXbMWexnC+khp4kg9tsPHenZYdbcDB62i4lq9kRg0LJ0egBG
LBGnx6hY28XtsJj/sWDsmAVJ/O708WJDGl7ojPi/DPQfkcbNVeVPsYoRzKc2rDpw6FeLS02UwpcC
fcxMGvcFWnNoQ6krDNPW7HuiPdAs7NpXeMCZhwh6Fpzogt+tek7I3ZmQisEcJDH/kFAmCzVt/2SB
JtlFWw/w4rQeOpoNZCDkhamJkWwtRk59LUVVJQV93cFFp5BcIvXEAPtMT39/Dw45Ib2Bvm7UfOg0
isuDvmQuXi40M5EdemUgH2a79C4fFkvYOi6p4jZQuEbsIKtvg29Nvq4aBk8XgZ2h8rm2SQSv/TD/
rxZZperiYUWQ4aB98kZIACo3rAvB8bMXplmFZS2gTHfQMlZWeSxXFB/cjZAX1zTxxWnwkuwxxRHd
vbSzOce3dOZG74/+7LJwWBSA0nlPbaUApBss+dzq0/SWPHpZpGZ3BHVomZb45wjy7yd7x1b4a1tm
Icq4sNVvsbn6gCvqelsgCy+TNQis9Ja8AFjgbonqEEm6+/wtfKKnfuWuYJVcyzmtyj8w7ld3Tqhn
K6sx3OIwAcOucNgZI28YHQbOuJzuF2oZdqzXm3uP2ECiTXD9fih7klPNY9dKNTN8f/HECgUPW1eg
GfdU85wDvDtBUZ9hXpS71xrO7K8GU3pwpSFLJPXOmsYBAvH8rAzKXolXMiQKa5GC/y6qQ7vuq6pP
Yj5BAFCMl9Cg8N4tQYwlR8qcvlUTdlPSCV8SRXNE8QM4G3lRbTM+AO6bl6h3gRSi5iL3va1xAwWn
9Xfg+m3G8A9xYGuN7bx/Mi1ZOW8efQ12kzxEMd2b2CGHywBA9pdyVKS5SPDC7O/0GTayYD0mv6bn
KxUttmjv79pP+8sVWi5yLx9iLJ0VzEK2F+sguKBfvxRWmnjuKfIv2GNOF/oZHdtpcg+tti82EE5I
D9is357gmQvhgDUW0soCLHqLPXo/24ZCgFNQ1cYpkv7aqm7oDN4JcjzUg6zEDIhb6gjh5HxNWhGH
Qj4ySOD8AuuwBhdOSXh51okR0HjUZvaB6oDPf+DP1bhgomujtEHPG1zPycJp9spSRb6AiTrzQxsA
hZjQH3thA2U//eEdWJhFOOPfXOKJYpJiDiAojGMY2OYsiNEf3EAVbPZ5xsLQbf3aYE6Ur5oqLece
xORrxDBk/IpwVEKTUdnBvfd4aRsTF6t8bLG3Yacy/s4bBnsHVezX5bP0M9uKYP35EKUd/P0Rm9i6
vO213sSNFS4s5MLD8JGKYB5Ez2vmf3RlHikK/9u8OpwDfbUFxEgODusE8lLDvCMWb1eBvqFk5j3C
YN+RHteaFTdI5tmiXy6EbL1Ngiwz+NCKKGXunbfKcxnQFaOPK8gCzF3sRfpPe2UmJVcnKM7NXpU+
65j7ZFVqQm5gH+mA/qAh2mo6FzYnEbzTmCxKPdPpj3fawAulCG85t6qfComLYSgSVDyYLQm0rdY2
vwLiwU2aBfI9qorZ1dLGT3bFTuxL/sVY+mfQB3TZLxImeMQaOdrYoJK29OKpFRDUeO/OkZimG0qt
xtgbEODBZ9R50UAVYdxl7YjXgkOeGiBIDl0m0L1Kswgx+C4/e4fU3tRzJg4I/w0/pgGG5cvWOCi8
XpeHNP0B4oOV9spRKzYtwF6EhxGb+PEZixMxOPlpV01BX9E3BAUpmx7VZbTK3av2BT4IbVElGV1f
T8mqSIv5wJ57prN0ucCB/ci4ZNmN55j3XrRFTNkeb/1O+xQcKOJ2H4tMLdTuewgX2Ev4cmVd9gyA
cj0nuyYQ0UwEIm+NQu0lH+Oc+HasK+oBgPtSO3ZcTw6ZJC/2s0F3bYVLIXyVhtSpLQ1+hlElfyuq
5DYj/GOfOrxQ7S6smM9PxT73o5Ay11bz34ziIHJCwPswwUeSD+cScwVOzzb63F91d2av6MFWPWwc
n4vvPlntmF2HMSv28ZgmUZmPU5SFSATgIGQQiFpaQA40IYHmu60r754RUhKYC/a3e1UCeVSUtbEU
fDD5FqjDFifuqN1kHgx5UI7sBeLIfE6cZ+4O32aXnxjBXfOGwQPDRxcYrcvig0oNYYwzsxcAHTpt
x8TFtZ9VR/ElDV24TfOUsSDqrReDQvW4oFRUB/grT6MONSSrIsDJeS7nf+DrEDQvOLwZO7i1anQ0
a39LgIb7czCRIDqB0a0JBfhz88wEPyBxOFQ591lSWuc2XE0+24JdJSuC6IdWGOwABoSHqXGjxczv
0ejUaTz/canPXDQaHC0NS47nj65yNwRiapEPE9AIPNjuImqy5sXpE8xD9Z7opwh3+iSoFIgAMADI
dgAyAOqnagbGZHl4mLuQtwwvP3QNQr73MO8isfosdJ+VoaLt4CTgXOwRMnljJBxNufD5GIMGil5F
gliCegHCSrkClRMy48v76ITictT0304NbeBJuLtsFAFJ5UvNv1bmuW0jo+SFuUzqoDcavunVhYHV
FYuwVsxEg6t4r2/FGS92+BJJfLdvWx1MJBJgrU0ZO6zu2jpKIPS1Qxh3rGPf+C88SsSCxVTunDMZ
i9XRJTja2VYTGXRhiI91yzMYvr4K9OVJGiVpkdZr6WU5nB7zJEDv9MRAIuvIUDJ64duv6m5NLf7U
twlJzx2d7EgrueuZZSWYLCOoMR5ODkg/LRlW0UFTmr5TJztjZFut9lk3eDgf2UzOtBkzBnxEMLO+
SIdbYRU4iEFGWZqVXN29S01rkyzHJVk5y8YNiLid1zqiOSS2mBjdOc02ie6HDFpq4VEIzKKEmgDf
EmvGTOurDfUJm1NeE/RH01RZyY8io+yZYRpRwLr/d+SnwUXzAp/s0uKVd/rcxZSspezHgvXbGyIU
sgfZ5ZYpUtZZKHeSyMuwk8NSot6fzTfDpdIowUvzRJbwlpjHm/ZJb2gDm3FtpJZmxPCVEE0i7n6W
qSPVNuPgH1Gb6fpWBLtMH2Ihaa5M4biuNiJA6GuP8d9WfzcB36jibaEuxID1OXlO1J1vRW57o8Lg
B/76EEyFTRwGJ9Y0T+rEABM06TIO/NQKRFE3PF8SLBJA2nsY2KQyF3LMAV7Z8UtiBOBw9bTYwy8D
+Um104YbfQiDN13g0+iLQ9w6edZVg7ppGRKLRKwpHjJztzHqaGIX01MzSXttuD9Px69HpdfhnJQX
0GlZaqH9FhNGT8f6Dxu/joiuUkbzgh95KBkRvQCJoifFR8Q6QDqzHmPLakxjXC0iMa7oP8j2hERB
9P7RbK/4iIgWpO5apVO7iO6u3MRNuqRxjv6uGqO4Q2i+1Xw+ivWJVJE+DqJff5Nj10OLWZfOHjwe
Xk4+H8/jKVNO+TanxhuNe2b8bLAFQ/ciSkCzb7IVk6uA9rs5vch7+OSebL8kFwK0C6BhXw1EVBEJ
YpqG6vqsB49hfCRoe97ZkwnwhnyYTI7IhO3h/tMqEF0RVy/0vMgFIl/XE2y++o4XY1XSOzxjYZgp
aXXIbvC7B6jJS1c7uiIH+oXDco2a4iPjP1cO52B+H/J45Z3acte6WkQXGI1U3RRdcnnk3eYDrsaF
zJepErYfTgPAEyi+kC8EnsPa8RdtTryfvZOOm9lpGJu/EaBlRzVulJytwG2le+tdRlB1ZiV9/TnP
Cnbl9Uk6AW5SBVsqQ314hdFRP4XY04/gVFyT0meYclIzRgq2oWFQ3mp9X+svrY+G8klpCjYLnyS7
fiDLQzfSEoTVHqihcBf3xOg0ZnXqI5/RU+KAY622IiOyvJdlClHiQDqFSZ7G7uhkPIivo/YbMcid
zaVY4xJdir+bG0JqSb44fB9s7pawWMNYiCD7X9e3GnHzigVCuWONn93ifFeFF82bvVUz0ojTUs1S
NS6S29zv08PHWJrgCsv7RRbPMXkCR4JRb6XcOAULAbdy2o/ygHr1cLKIfXclvSnurauNhF1d3yno
fN437apklbzXOR7asYucuFY4KncdMtf+9uclORARXYSJgj6Yu/TFGzxqsVM8mpAtwvwRhYifWtnD
0W4NCwi9yCOAcwizc2bbe4vob/yOw/NJCkww+mD4j82z3k7mJA6igsEHO9Sm7dUOMV7CUM0N7VYr
i0ycZV/EgWGPmud9NBqWKENgpb3YzjNW+aMq1vNkM2VVoGUoyZJIXUytmVRduQ/tJaav9/9x1g48
mMw8JG2/YlsUM3Se1k3KMcLXWEXeP7s7+bg21ORIYXHC1O9X++z2hEnPam1Cjf6g2aYDIazNGruR
7byGOcLOsxPuxJ6TvYjJbNPJQFR8nPDEDX8Y5sfluJj7AXH68sPTJ6g8R3jaYfkNNl8N8VTSVKVA
X+qEubaQhgSGrUamcKwjRIjJiNy2YE9bIuxdhn79njQV9SdtDUHSPVOPUbneyUsNjBbB5Aga7D17
n6GzOepKu/BxtzsVl7TWe4ZjbbpJgp8d7gzuV9ge5zji1e9jTs2MQ4SRYjoj/OkTqAj/4K6wWTcn
bW8+rjF4v392126nX57x71K4op/YfK9PPs/jEApkftJhbpv4/+lQlQQpYAH9WRV+8y9nCcyfBycJ
VPiIPeIR98ZmsaVTItmU4K4Lzjpn6SY3g/C+ndOOjySVB4SRTicYx1o7yhMWiYJQUXpIy+laSUa8
9qyalqqXr7L5BhB1HCBJg52sKPhPSB7/i9+HllBjQilJXTC6WqmkkRRcfLkWQ1wDe2cZzEoxMJPR
79JmTXOfQiKA4McbHUsUdZcIGsSgMBdmYmGxpmJ8pxuEesxl9Tlk0rzhMnw07y1IYQgypa3BKt3u
ipPOw9NHTfl9OBwJmmA+ZntpVgmHRe0R8g3uXzUluwzRZrm/e49NONolqdfX2Q07ADYKwz/kcYv7
6+h/drQFKpBwi/RLtGLDjx8iHxRnoGmx0IPXp2CtbUU592bBp4q5qr2gTzrsn44Xm5LgYiwSThyc
jCqe6cyIgwvueatFIRT3VJ6lQwnHtRSDg0UMkWLDwRHFZ8bSy/aCjz9PBMxgs8NMP8dplxw83src
80jrGZ2DX2CozlLCAnapT81eznRWg2+p5BVwPiNuzv2yXDX9842biQ5fi/f/ryh22NGdq+hk0AZl
pVIkAc6ybVqElOPjbFASXyt2ZHKB3phfT3GLUbssSQZl7g4NZTf+tNoUIaL3utpdaAtGoOkf+bN8
ziVto6O3LHAxBarg1WSyMmS2S15IkxwHmOrZi+8TEy170MwZZIL+d5xpOqOd2UecxUFQtv7euaKZ
qRAvkvEjE5qUcKfkH7KFKUSKtU8n3U4Zk45cf5FkdsLy2uXj0+m2GmX0eX/6M9G9YvdNPc5ZPDV+
3giS6SENsOm4RbHYoaWVHKqZoES2h+yhF1/5QrZ/ARJI0R9207FSQ/i/n+TbNLm7x+XoLznZDMEr
CVMCggj4vK8+D4YZiJY4eQNA0iws9G6caKOTBEe1unWsKMfgm5zEUyK709VqgRdxk5zYWrc7mQAa
iqW4XT9t6XsK0JLUzt8boWjK3HzuUXBgf8FoQ4rUDGuxY62Bw1QGNokKBh+OFv3SUsAxkZd/Rhm/
Wn9p6BHedIjl/kis54mrdCseaYLtbk7QyVgBaYL4On5Ki9g+5RVgrR4PwtNgSWfaq0V0MUSzM5JR
E+eytkv7U1hspkFG/rNWtjO8OQGj8VVHhuI4P/lJVtJfGwC7/ViLAOvF8yVyhG+PKwRpkz0dNbGZ
NSurOUuPwDzH9z5ohIzMMxvyrxiXZtuTML/KKeffQnKyZoBkFHE5Dlq//lmSBgD5XY7oEmfpsvhM
1RJqDyHOz7/kmmHDaFw7oHszguEeI5B5CmJi1/iR0OqhxYG74eofWd90i7Dd6l1A15gm4N+Hd3k/
FEgMNtN0xXPpWE/zyD3QMJFa0g9Dg7cpMhBG+Cqh7dXu/m/Cu8LT6o7j171j4uHdW29YWwqpZT/w
sGqGKTJDiaumsMvAQ3lxYWRtW3+aQAnvn4MexeuVKy9XaKJkIeBCGumsmnCot4fvNxZLii2Li7vE
JIqUvyUzOwYX89LUwG9uZ7LMPKLlVIXXdxQDeXLyk1ZMmrrb9lzR1YSE+/RjsNiHDgfNEBSEdIf4
q3EBZtmrd1Kz9s3L5XvZjDfKbPXQhNcCJ82ftStfDmZFC7WqwC1Bjr4kSgwN8jBTNS6DeqwlL3GB
oyIH4mbNYTyx6vtXGDlYQ4xgpLJr39WKtQk5uEDmgXR+XlacCwP8LYfiSS7fvLVVB8j2D/ABf1Tm
/ZLHRBjbw3xUXiHmiwLkAVsY6HZQJBlxcOxZiCUFouvKlbiti2xtkjJP++cg6GaBI9KsLPTklUHL
I8dnOKKmZwefSlMWra58YH+wO+Y50ew+oXyNvoGTJmCpJwWGmeugq3eFUuHZFe6GuWL289bvCctW
jPBuOfRsDbO8UTIZld2zmyRT8FNdtiURMdxHvV9D2epVh4AGCNnr0yydszV47ZvGgDYWxsH+kE/v
utY3LE4Z0ekzKtY8RGNAT0eIQhhPQ+KTWQWF6AugGSKXCAdRP4kAK2eVLjjj7mg6gw9NdOpjNtd3
P6WAU9Q/xSQB4cYc+7oN6WUTCDh2W01M8opW5VTL8jvjvFzHwRc6RFZ5nhwD1BaBk13rg3T4JZJR
NG4pvuYMca3L7MuoOjGi+7AO4dYNfcqPjfZ5HbibYC9MfL1dmfspWmiEgFLk4T7vmtn4X6iUDnJH
lscaYLRebx51/shlq5AMaSqPShjQrWCsxBtXZ9Jne5Ij5RnixUfF4oRsb+dXTIPtafQvgFSRs86y
m6ycC50Cd86PPnzs3ZmM0ALlQCFGq8w2uSSrRnA/3bAQFa5vXYZeQNoFj1C25EndZGcKUzjTu2mZ
NneA3J8hwJfGFjBbHkbWBqkPtiR7umzcdUNy1of5SwK2r4arePXN7qWkkvwsnWWAnV2v+F27sJtx
xkN1Uil9rrWuW1wq2W1rozjdjD2H7Hjqes/d1DQcZLuESfBHf+1IboaXVY7Sgn1MQvbMGvl5T/Rm
l9Nzjd5UEf+lGg/n2HMstv2oBgg+JG7dArXzIKeB3ZXrSqhw1uRUalcCFbmp/dX75IAWz1PN+G+k
LTZvNrxEAroqnWHd1xEkMovlzGUG3+SbZL2ZR4X4QEhwCZU0JMHnhV6LyD4U9tHaAhcBPMbkIa1D
aieo/KO9YQLhPHPA/6Tb71oSZw6YcndAt9PQsjzmlV5touOzuRPJeiQJGUhgZe/vp43vYwvSZT1F
CuhEacBg9u9cias0c/WV4Kt+m6ZeFH6+cZZuq1Hp91dcplb1F5f7kbRn1Y9p2c4OeU8bVfcvlfBA
mwokoJx8j5Rv19CH4WzZpBZbI7LXLA9cxBnN1kpyrgcBiCr/8EC6rVnrJe/1cEwjkgVhfQljRu65
I1GsUGFXqQPgvi4Z0TTNtG9JX3wDGXoJk9vj7/zpA3qbkrFjsGBym/vw3FmWRJtePa/slc9KqQQJ
/HvhRN6sEepedHHViD2ZayIMBVwsfxv5VuYLWssWd3vWkGR0AZ2OWLx85OpY+c/Y0She/YEHDOdp
JUMArP8dt9gdlvbTgI6y2V4D/UJhvj175di2QqiYg9jRg6wPCQEFdiDI9OftMkRFOXgYSdE6yzF+
68CP5tegxoOnKjWz/qBZT/hNvfeYJBjeZN4Rw4xxAjnbjV0y7DOBachA/TjBb8EGc8jZ3Q9qwlAm
ExAGNdryRro4OUVzt6pLh+2+msk9DRZfX30pbw4ZBu18DNd/FwBr5ZGRvwEDzWi/zv6dlT/XnAMd
EQwx2P3Kb1XbJD7K5GcMZ2ZRaGghHmhANtJEIYqK0dEEES85x4iaBqo3IJdQQxkpIvO+4624KzFl
uGEuxBh0M7ebxRhL2yw5vZzte7PsSOyFWVzRJqHp4QNeJdE4XViT9PIU9iLLwlN34WynqPj5uCIf
nrUOVlaLIE6FF0bQ8vMxBQotTnSfUes/feD2n0tQkHzTC7W5FIOXBtejQzFxDW8j5gKJiu8+YybB
RhGx0STFro+MnGdKPmx+pJsqQCmFNFUcxGZ7ny6Y3k54YlLX5R28CwQtI5QAR07rQSXnG61t5ea3
ZTu0nd11GSKDvmmJt+OAQtu8qiqcR7EepXum27unBPDfFUHJNI4UqrS9V2pxX2f94QW+u36Zqsrr
y30cUifd7PjfEJKovsFCHgTFWYoqpX7cqSxgmcOAlFTZzhN5eIzgqc1llnlJYFzUeZVmz6mxd56Q
pmW6uPw/iWHo+RC9cLdZ2OfojZsDreRMZqyld2Ho+2YzCaXEB1yA6BqDan9PS80NV4tq/wICUieC
BeQkkJ0T+yHHroEdJUnocMaoj1jS2xPYaTborBVld8ib3+j8RyATjtfkyJBfC0iPlg05yK7ZtFM4
Ck8EdzGB0sNGwRt4qGhUI7rt5AKwteeq/EFp1Rpbi3BM4UoI+zDOedYLO8dqNViuEKqtwq/NPtpt
fn0EQVbJQaFwFAFCpUqoPSnuoBAAn4I08+GlqGvOVNjMk6b946lx4yQC1m12qzSwCmrG2BeDOQOD
a0bDHmQuq7T1y2230a20wz2BD7gE/AGXsZouSHHnjD8uQEzjXpb2P7JcL4xL+NxTWNWnRkeagCoM
vgi52RLZdyD2iyGsjXWVZjYfitsu6AX7I24UmD6Dw1UYQXWzlg6/MbEqWJzNWWam5uMLNueeu9hB
+i+PT3yQJKwCxlXpz7o5ifQN1ezNq7CenMt3G2A7WMO9Lw/Pc/0jrXKbw4ueA323N5z5oMDKQMgU
9KktfczZshr0+4zP/NkMwT/LqieuhuVdL2f4yVLCFzNAh2Rq368txoBNTnsYinyg4Fvjz2H/T8DK
7NeCyfcst6tvCmfcUDx1LKazoYU+KtpHn3CL67wa3YxfZAYWxUCD40DvZZied2gq3KLRmv64SWgR
3+GAskRIcAyRpzqCfHpYwLXao5kr1w23cNNWIneeAOnfUAGhqMyB4v9LfUSjr4wUZUbInN1Lv6Zh
xQaTY2Sekk6wojT8k8kz1ZWeNuLWwmqQKOAR1RQmyRFDQbfkfgvYOV38DpSoRGhMrnGmyvLIwTTj
3zW95jRvZRO+L7qmckY6CTlp8HaKbrG88g8irk9UMcwOEWPps30Le1UZDXAe6Dzb+4IR/sOKDjfr
OxkrHBzDMa4ETWvHv+rYsNTMMa+X6tDOwXGnU/51hNonxFlbMZ2MpeQ9dUJ4YSoKK1oPrQdmcWAM
Cylxx4XzTDqwe9zQBKNg4m7KJ8fOrBzjpaI8z+j6nEV6lif06YYl38XW7A8v1uHcXKJFwIuuATfk
lPEB5A/8sNhTiRrjDPL9p0+LC5TVZ8XRUWVtNwFpXdcOyEJvOqDs913dag1HDYFNBds6pdex0igQ
cDMiGdAyHYW9Gr8vniYSZPaYDcbv1zNo9oZ770H+wabY/PRHmcXXb7TtPes1sjsD8ook3SkOF+hk
Hns7yl+6sdspoG6KSPq3052FZcmGZdUdCtVTEabFmOG3dS7UoNXl7BoKBdZkdO+DxMB9e+nPMjkF
u7nn0TTm9j5sM3kXbYiXAkMWxZVMi+6hzXNdFOVT4kM/+BgB0a6bXiwCTzL/hPqwiUqhri9lCLyN
62uywRNtBu/1XVXGowZ5tRnerKpAA2/qCVQgiNfFnOeo4VhAzfrFfU45JiX/k9NsFYerGT/1m44M
Ia96vZBma7e4hisllP9JIeiqr5waIuP6eYOnBfdpqY/4L9yD3CdijsUxnSHziZg6Jq81L2ZoI5bY
elROepUiQKjKrZ7/i60kcZrnGBXtGXbFU6Egxs6GSFG07JmER5z6wXVLFyNsfvSIBuuI1jFTRarC
COcGK+1upO3T75gS7jCuwDY0hpqfcRctLQzL4voUQHmbwM/nKuBqBUJ0a8CxpXpz1DyMDyuvz2ct
cFPJk9T5sKF+MVT+mYolwwqEwookqZOVpophWCrjAMj0DOxWbMSDKtlSDyYeVYAx86I1KTTsPdGb
p4SK9Csa1/KwovgUEBYoSUvoxptDLim5cJ5jc1mAi+5+tqj1lI+cyrJ5v0E6bvprGQ988fSjdBWV
q2OqXHFrNCboCdclJpiQykIbsV44u8gvb8sKd5dtQ89HQPLS9FXqd//mmuPVJClmEaWHaBwwkYcX
aHWtLKCxiCa/MFxRIHQABWOE44D7XmUdLXZ/cR0cqSFesLS2UAJVu8R/IG4XOWDifMZWNcURhDoi
IYLTbmuZI461jEZrpeNNBjss1mYn4RKtVTFoRtGFGsVPUyJLZpHzdRkPrFfnBMJKqAwzrQW5q84o
pkDaoB7iJmkSn+7Z6kwqvTIE+ovOWgbF/9ar8uv1cyr2d+s1gHDvW61sNVJYunLjGvEVX6GxiY6C
H637TBjQUAg09CReNd17mqqkRaPxqJ57wX+JmNWivJm+VkeInSoiB0+CydsbsCI16DAB+5yBz7r0
QPxVGxGDLZYUSu5em8c/Vr0GijKy4LoZD0NX4oh5WFBYgxGwyjmo0x8eTXEtjZLK0QyJYjjq8RbD
UcCCLYlyK0hu1rt1OnxyIuv9XHkkiqLNRyyKOHobGn/EFrZ7Kwman4oL9+Vk06WlVJEEcp9jCIRx
BNesZbjI1SomB+Xz37QhhcK1TIEuNRiDEc4n0p9hq77QLTESkIZ6lEQmQd7/1veu7dmJGvCUapMC
7xb6MP5zjkgVbFAHSBy/70EONqiPFrDIiVRIZBt+dK4VsV4JN81ZoaPRcKtMLTnHa4ESTTg1XPeo
UqkOu58QbL+ha6m7sA0s3IWEFh+LFm34EOmbnacKIB4lSLewG/np+jpJBvrMRlLam/9wjm6iemrn
De0/mBGqKCBde0uCMDaWwtjKhZ/wCj+m+8hH0Qh4aEMWBqTC6tLrvcMOZp6qUCg425ZgdvErgGwt
CoEIMsHFoakYHwh/8bWD6MpoCdiyvnd3BaFoQOFZhZZrx19mRqxiUJVTVel0dwuCWVYZ5DaYVk5G
JqQMV/IeD2c5rjJG53FSPc3UcCSPQ0516pPRq83b7geN+IqqZl2fimRAJPBpnvrj/K/EKL8PFPN6
vXPz4WZ3/rnZ/HiGnhgSCrp6i51llBiNskZslQrfXjU1rPSdwRrbIK/D+urcOpgTnR+u4bHVkV1F
NDyWJJFq2CcKxSgOBUk1DHwFc+FG98YvmMSAT0e6Pw/BoIuL6A//zFMM8UDF2+CKLtRQJc/nDLdn
hdg+0ZS6u347uWeh0ZiOUxjE6K66i3MmcDCTQm2pGFELItKO6PKDbDuia6h9SL//LhdAv0+U/dJI
rCQL8qa27j2Mlr6pUtYSl83KEYoJzITLiHsMHZNi8Ib7Ma4H5HkrMOtKkhbbG4S+840Bs+1fk6hE
ykbL95G/xmYkJQELTwuujy59TEBK+osc2fvG9LKnfC7a55SkBh1e9wOW4fbxOnbFoSUgoF1pz7pG
1P6qbpX53h9M7wOs2f+crWVsrpN3txeFCbAewT68FQMAapqbUBZ1ASsRALqwlsIvb2MvtNf+JwUr
7t4kLqhQPUmHtdg8dWrLBxdXjx3BFON4dxz2oAXUFI0n8LTDgi3L75dPFWZaO64Mo3c/Bv8GBCNN
iQjnbheCgAoZmLn2J090L7XuthEhFbwRwhM95G5C95WgpTONPZ+nNGt+NwlpGwO/3B7xWeqZRD/A
ySvBIsnZ35YpnStjXza25BwU5m8ZlQUDbz1OjVHbmlUEk5SCEBWkf5IK0Om6NYvmaOtinsrnAKtX
qRPNFibp4ipDJbRMKb11emtCwABJ7wiON3+vsXTmUX9ngE9kFWydVe64ovUTqrTS3DJW/5KFfugB
N59Tli4orT1jWxRZpGIagTB0gYKBf4Z3S90t9XHlCckRotG2s4z181xvCo/gskzEG28JlRmrWMNL
jQ6PkWhTPtNOSws95r7oz8i2OCAtYg6PfsKg6gqZIyuZ4x0M0bYqgpiNeeZ9TM8IFcOg45mmH80j
4FYAm6G0NiFRkKfexslf8+x2Pgn8rIweqseE/RYwrdnRcRFTALNKb4vs71zrxnHauS05OmsvEdFB
NFSKrUArpGj0w+E7mgffEO0y+eHPe/Z+ykcKV+0L4jgw+E97HOwMpi+2wD9qZ0i3gPP80LoRT4K1
yG7hxsM8Qp1fXDT6BNq9DwY9xW7RhvRiQyf/sAp0gFS//IZG6oI+23oVr/TFWB2rvB+74S/PsTsF
yH6V9hpQ9CX6IIrgSTIaUhtZrM0ktUiDnEI14Y1W/7xXjJ9rY0e7f8ZST5zyZTktpkRkdwVCMNYH
OG/WSXSeK7q5MTw7d0L7pQ+hrgOEVp9aIThwk6ki8xkp2SHlszTN7vFL9u90lfopsp8c6cUhI4Xj
e3nN1XSu2Udg/fKvJGPhPb3faBUr0xyr2d/FosVFNPBHL4OUpM5oGEg9Kjfadvk40QQGUxDgeu+3
PsotXrhwJgXwwDzs8Uuspq/e6LyC2IPyygGdvH2D+cH+NWTqgoXoNXmvP5dj71vtnTGRTVgDWp8q
XnhjGgD0Cq2mCffmazrN0AwtfNGWpPG964Rk4TOOhygVJbaW5BhHlcCf2PgNzd+wxuPUSomBziBH
7Ww336BGB3TcliJsYucjxt6T51x8FIvaupJc8MSAyDkZhLJbsvypAgpmZy3CcGAS3Yu+qkLneyKs
RJ6/WaPKXja7Mex7YitB8uDlv6UfUxWzDY5tVKZnxO7hRd7qLtGMwqT9GgQ2DQaYcx/kZin12r88
ovLKObHEUASG6FE7/pc7o5Tb8D95yIp7Vg0bkojNOTZ8tLM8azg8UvjJe39aLc2TRpvt0GOU96tO
oJenUy1NmbHd0cQ5X4I2L7zN36/wkJF827J4Sa3yUZODZssqNxAEdwVSxR9syPiEwU4EZENcCsan
Y+HxbZs2DVE2Ky78UObnBvWo0q4aABfnOsHJXNHAwsS0RQDuEvHiuf9kAk4wiTENqQU6mmXMbAL5
5OUiWxumEyOYweo7XUymproZYxkzfDsFqdHNPv6gt1Al66nxh2eULdAoBJyaFo6dUW3EKZOSxkF6
uZ/xtzos3RWHkbUPLnPSKO4tnZp2BiuWkgNNme6THSrbkvyP+w5EkdpneSYohL9IcUipyo20CfGT
+yPtWjGKuQjipvJdCHaIsO7uxTORjCfKX/FBBafqW2YKYsXUV5mt6KURzmhDYAK2ePKiEEJvg56Z
/iQkmwKXsEHmlfsUyPecqqYGKlQPAqFic5XxLA4jIXP433cc/T3vag8lLEUmgqTEkGMm85DODRL1
8EZ8nj1caAPj6UjJLCHXLobYS3ghDThYuojI2JHMhHLuqsixC/CBl5B2lk3CWOlJF9eggMN1ALWm
FJwk5ORn2ZdC/J+VHC4NGUmFCH7IB0rBB3+fmJgiUd/Ciee9KnUNOxrq9JXyTb/wEpdraePJfJWr
E2j5aSzvtOsGI6dKo+rV9omhHUdoD1oiNbPX/8NpDWu/og9S04lKEeQzeQ6vVqrE+WCH6diBNPoJ
VUp1ms6lV5QDorJJfMQkUMj/a/EOPlRG7zpbYO5/jg1YpAb8CocigO8V8QZjDCbELxZS0VJteQP9
mpjXVbuDnbuweMU0m+mJAzKZzTcU8WJL+PL+K9Cuo5eSkGhOyyLRWdrBau6gth7dnJipOHjyyFi7
QZtVZDesTdSHMmu7Q8m4jGhdsbCFcxgBjRpKBOKxmObEZHcPqg5bBUsqXrfp7BWuf/0wJ/DgF0rb
MBAdvGAXLnvS4crCJAXjQgqaFoUTxkYbDJR95Uhh0MBde40MrKYbsuJMPhhnRiXjRc+mfu7EI+gs
xrjHkvlH7BeAXz9zn6VmkbuaGcCAk2W868giDCUOIw5sb/2VjHzkogatkXSHpDhLTj1VfO9WJmnd
+hzaNDZGXApRmlRJPR/dIb4ZhW/2IyV2TGJCQyW1kRfQgOXxLTGY5gL0+4Y8z8QNmwgFugf2PRt4
AU1GTElSMHnROB9VMv6CM6MlAvLBCHDPyAca6CMT6dacJp/xrzKhN85b0wWMju8OuodjqKpmzJUB
RDNtAEk6XLB/l6LZkytK6ePIEAXb7Bb9BrYjjr/qzkO7rOvE4FMtKZITEiM7tzPKU7/HwQ++YkTa
TP4T9GZLAF/qfU12jMS3Hi7fuOeA2D3YDimAn/py7BnI6QwhGpotj/+yM7XvMRf479bZRXRleHC4
gfEjowjVCmH4O1XELPbmJ8mBT0qIHl4kH887nyd2448fb8HkIaQgtQ6kjSDj5NCpCQhlcskiwPOg
fA97/cqOcoJQTRzNjE57s9IdEjg34fGqVd+4SuAXV2FPsVbpc1IbVJKYy3LEHtaDWbBWHyYNruV4
YaSy9S6tHKN66poRV8dn3TnhhX+qhnyuEXy5tBfaIBWXVChu241+jDIzpnbDlMcoDh8j578FVdMz
ql4yItONw9x+5VQJFhEJnZZ0GlQSe/tnRabLqAlqx/CeD6hLVu97tlievWyVswgB3wlfg7Jjjj7c
El9ZYq/+HaGmAltRtYiork2Sqt+KmfPupYM9EQjxFv3QY7dA/jNxWNHwAlO4TBuh2dY65SDsJFy6
mt5Lgd9oscXYjSuXiekKxG3j/VnZ7/NkthLbHrB03eOAwASE0xQOKuzW3F+5jQKTTrLdupr37BVC
MpHzSE/i4FTW57uj//Q/xvlZPw9Bl+whz9oK79VRLHp2nKVFDKLI1vclEuSQgHzUNa2h5Dpc0mSm
U/s62ToZNnw0KKPRdx9GqDoP7X2uMxSwGmN9zGIPD/HSxw8RDJGgjDFrHcxjAsArJB7epwrrkCGZ
J/6DnXP8UsPgNwIgK5RJwYMlBUeSIIM2wDVfWMaSIA5DmSQLsgFWQZ0epufuiUe/GzROySs4+IV2
BhCo+VeSb6ankhE+j+pl7vBoFRXGw8Q3vq2hzlRUetuB0q2ekJGtzT6UKnsavi1eJiO8txp38OaU
qmyOC/meR9eow+OcchFCdgbbZjCTfqVv8xCx5cU+fMuw1DxvLIFGw+JBh3xtBqSVqlgFkbQXMvp+
pSySnUPXX4KtEmjc9Q/2UMVbT6hSBgvUWIFSsemmRjJb/lI1RkAXOLZpQ4+WMbhcCqLwqJZWqlcb
qoQc4qp9tpVNe1v3sBfTRsDNbSOtaLbKRwwQYAtLN2VxkWqx6nc+9T3paXeueqmuh5luy/QujyK4
2gW1JKkpqbJ8e2I+xoP5W/skHsKuuVQMnyzPIIurOEs3/BhQnc2CTneYKmnU2TIP9nMbeRlts4OI
fvLGEeHFKPqwiFd5wJBrxR3GeaGncx0m0T/nA/UFBaWLzEddIfHZyY4W2u1BsY3VWsxP9kMT4Tgy
3gODXwKYk4pQy63gk28yeNlMJRU1aP90kAtZcII59wXAi70FCKfSiCMJys6GLahNBg/uAqL92wSq
FDfPqdegekUL16TAl4OLh5MuZs8UmcH1PaArMrCr4AM972JV7EJdmkgPkjnVMDjijyQcClO/sqfQ
ySrpSwhlbffPwTE0HrH17wjOLlGfqYGdUhW1vROzd7CQV2SIiMs0dEPIlwBB2ALyoJRpY1PT7VpN
vR6soxdo36fVlbyFYUV0pVQAaeTeVIhHRctYTTnfn8+qkknpFhtKs2tBTC3RUHNJ16H8hl6zCcn6
PFOkifGw3K9luvz4D94IKMd6JzppovULhMdRTBDx09vFaJWUN63Jnn6gsWv7eQgiB1CN/CMYPg2G
8mdfWGk8SBoeWpEFRAXf7tsABhGcpmCzrh1tzUoBROiPJl7EFIPpT1gTr6JQVn2kEKGVPqhrAVwn
QA/JcA2SPalPA0KcFhqaCxXHQtL947zE1QcxSN3TFYyWtvNkfq5t0OUntKvOfTdhxOHxuQNca1uy
QViVyxl34OVq//1w8LHeS+A3o+arX2en1UmsxadnwrnwJqnuYQTh8i3jUGmSGRbEb+fUJ4NZ6MbH
QfS5AXA9Xm4+VtTHMqbCRKmKM2ljE88NlWQttQNAbmgMwFdDa/0SyrbhHwdmgRbHiTLYIbJIkdSZ
y43HUJWJuQQCv7ToCs4/r618rZO8p0fc+Dx+w66LrWTrfhxRWCRNDZu6QBEOOWVkDvIDI6Y6zNq/
1mfXYKkPK/yDw7ww5GuHVIdnN0SzyCHPSI+U9b7MnYeyr+6MRhuo7TfSzYXKlgClIz0HdrS2llEd
/7/8qJhwmnR13OflGO86dtGrnbvyvnOxKz78epMh+pCGp5DTpZO/uwqmYVl1la2oC17fdeEb9beW
MqTelKoJ+JiRWH7CwWAi6C6+hGzEiwok2epjTzogbLav8EsBWc6YQYueWLNinXoVMOoNHxF6prO4
O8RYPbHaHK/GZJ+sNHKCakHiRkl8sGUkRZkpc72unL1oTXkNN3xFZB5ylEazlCILvlF4snDiLpGl
TrDEypyRhK3f0ZABh3s1S4/FzGQWn5Cn26GKt1kK9NEE/4NZ32XQNqfGwwI+QSQlenZpWWTwee9/
Uc+xkBL5tQVfhS7xBZTqKDL1i3UE9j4VxLPxPKPZstQPie0SmYDcCjn9sYTJjAZM25OdnRaxb7/D
3mHvn+Yqf7YWU2zaBp9LxR2U3Qbi8tcYpv0+G8KyqSrkuKrOb7w1MjMdZSZDMPhEI3NtONusq5xt
FD2BZaSRcAdDmag6K3Rc7/O9uRWsXTyXecu5eT1Bc4vEKxetpx3SRmXf/hIu7X2zUU3ABgtIldqd
X4+YLX+KGslDjz/MPO60YxKnJuz/DNeaZY7iL0m+E6D+XyYAWdQe0R8azBVyQMpVD5LnVN8PWp34
97bfNVuZV3edh5Mby271AlI/YXayuEoyPu4qTd/C5d+cGVS5Hd/WSDE01dq+2lHyK98T9txJa7oS
u6B+dgN5tY451mVeP5+j8GwzPOUfPqr/hZdpW8jXgxlzuPA6v7dn+b9O4TyKhxyDNm35GQWF7YCN
Wx908OcImQMRI5F+MgcMcm2s7dGY38gg0bqYA1ygwkXkWaAxTMPT4i344MsHUuWVIk9jTBIhDRkJ
6VVlv4hS+acTVjxlfEIYYwJc/XOh6gGp7DNsUt/gHwVGxJy/Opc21s6B2rr1ZRLuQIEkfOmbi4th
PP33RIBHTQEatCQN2prBQDg8XeNDZLf/yvx2bP9w3dV7WsA2k1YpXql3NsFHmo6kWdrZJsw9I/L3
ziqQ5ndpq5969xqvm6Xc+Wn3sIWKhqXol97drVq96HzCrsM7MS8+jpsFwXmWixokrQPqfxd1A6+H
dh1mwAZeIBasl3BiNLoh5u0Q5ZsCS2fXrtc9PcK4cjXuCaxhBwbFptjHZF7cwbTqSY1zvkb5/V32
EadAZFJtzju3SqZa2I0AMTu+CoCzq8pU+TOtRMdpGNrzdSjp7kmJlZx/ZEbUpFZSIxj6Z1qRiRsr
5WjARasrl0MvmBQR+cZWbQXGbiLiO3coeeMYTWgDHBlVHdmqhSGw5lr/2AaRgHUduF1LXWdoTB5k
XUyb8ZZrsTYsm7a2k7pt2OoZd5GUYRExB/sQ8Gnr2W9y9ArfY1RpOnI47XGya/buTU23jRHFJdUL
2N8ewtBQf2PnK1XeVcLmq57fLJxeHxzUK6Rfd/eYrOtYJL8/MBNFuxE9HQ12M3Xou4McfovgYkwW
LxCDV6jbaM/Nq/btk4gSXJAf2i9XAnD8GnF5O6jcoHQwOApox0agTvNYxC5kaJGbupC+ixQV3kjo
9dt6xcrTL/RdPI/7mfT6pxf8TZwBxkj9HyAHwuvaPDDS7U+bRULA7V+wAH8+uGA4uENb6Womw5QI
NZQ0Pdj0K48R/44JiE9urZ6HOH46ST1D9wXLoz4ixhhZwfsTs9I4EMZhsakUXqv6U4u96yL/ThPj
tqTfbGCMRgLBCfrIlVr8/+/r83DcyC2ceezD/pQqFShXTKwVuXhM0QbVmQwm9hmzZEDJFHesv6b9
QPwKCegQglCGshfrWw8rIHrUWkKXGZxjUPYeyWUdcZKGC3D6YljI15YNgHPUNw8lje4S42DHUhrW
RkN3JBcc5O49V9ClwFu/+yZRKmgBuLVVMeUcDq9FS67aaUUdVtn9KMwCEZHt6HmhBMa2A1qtaY5x
vIa+HPs0yMrlyr8jMGsn8F2e1sXmpWLOxgZy3GyyLV3NjGmEP+ynGxt54XrDhb6mSYxZKKMRz95F
ojuRhQgxKA/2CGUp46Tc6fi+3wJQoRw3CNroCCW4GwY1USoFq+InimV8L2NYMH/RO1+NGam+RHDg
7PMpiB3aHNsq69llnhqP8nb/dgfV3ITG4KWNokq04VxpvzBZtxa0BbCPuwpYXbzaEJEXtAnzoyl2
jOzNfDDCRKs21ednR7o4K48sj0H0L9o87qnHEIlDqY5Pcl+JqM2W9NDLpDbEjAvLkMikex3XmvAd
enS7g6zRRu8aLsVbzk+4LZ/B5oia27qHEI+FSblSMUCNcUt4BS+YMs68levtJoO/xj8FCZXya9C9
IKU5WBs00eBnR7Lr11dnfuvHrTQ02fOoqoKqIKlzzYUn7W9GrtNlgmNeMsJ3Jj1mLIMMYGqIqvMe
8HxFzpWQdlRShh20bz1h/x9Me5EZfR33IPv6qHT0oK5Y7WrQMRtOT2oP0rk118p+j97LnO5hjpuB
GkLCy/EWVAh3oEBHP0S3/iOk6wL1KiNoG+JMOKzBt24WYRga9aimysKRKiQfAvvxv9oHANPiz1RZ
cGnwyIm/t0ozPSsR1q9wHfJeq1vjySIXrCRI5bYMBQP+VjbfMvTBEOewJJUKucZeA2AB/ZdgVo+5
nYqNZ/Ni5kxtnuQ4eeBWB7sdt0nV6ywL3dQ2mZ6wMoTBWgtJ8CEIbrnp8D+Nq25nS14gO0Q9mPs+
t+ZDrWr4OMzSU6D6Y+kZo5EukC6wKbVhWIk82ohPUhGYsX2v8EH2Vzk9wijSJRXSSBAEK76APk+g
h11ynjGExhecGIJ6Ds/6gbsqMD1VaYPRIPcUv85yFWp0eYbpMm1iVp0m5WPtuYo+InuNCsUID31Z
Q/oQsG9/OtwReDoXDkVq/9xyCk3fef+aoIPpVi35CTeAIQifgag+lJ8XIY8U9++iNRx+F+rJ6HEG
/oUNnsoshejXl4bB9wJvXAxGurCJ4Zi5W/VOqqweNTFuhRXYGdh4HbiMxYleocpLhndvMZatOAzW
PhT2cv+O+Rl7vi43akJxCDv6CpdvyPdgKCpGq/BQ4TppybwfGgOmtC5Xp3y/D0Wzz8C+UvbdKEzV
HQ53T+0ip2vQAak450gJVV3iutC0BsONZO9fzDNz3b2sw3wfcSi8p1ZT+KIY4X4wnSGIkSXHXOe+
aLE+pT/kYbq+8QeGwxyphgppNtXSBZxw8GRaVkEaoA/HsFONQIJB3qcY9WmU1kGSmzgQBPtpOx1q
6KHmHKl4m+kUEHmbjo9CAYLGLsBOWbrDVZpVBcaKg/1fGEcbQP2pA0FH/j+5Ma1uUzjcp467osK3
FLMRuhnCAwu87H6KbUqObTEiYwTvLf+aRh9xl8F8UVC0I+al14bNC6yijLinMFQuRZSEJyjA+8zt
X7igY1ryTpqQtOWp/ShzPYImdFU5SgGmmSV9/PlRsNct4B0qtiwTnKJGCgoJd5USAZi8fIziYLB/
Fd70RqehNdoVh1+y0BSoMjMPlOFVRWNnyPyX1oMqAHZfGm046ITlz2JH0AmrQjzkLd+qGfeNJhcd
5/4IrNvJlgSAt1PKllSciZc2PUFZ3hqnlyga+oPXfvKtf7jgbyhLoVP60w+fPzH8RP1zp8fceEW1
f/vKQeVLjtGIZ8u7K1S7O7mZi4EpIbJa5qGiRsIwGIaUQR+/ew1JXAjMVn3DWQAZ9y4LOHjS6wxE
3DCaRTnddYtkYLbq0OTcqhGhmT+liM1Qk4hwBeYS3kaAc70+bmNo8KBPWg3RDkR3HbGf8p1/e4zG
8rBnzHy7nFdyITOthWI9m//N86JVN0jvyElOth5BAxwwFVzhga49pZEJcvSg2YwMBNUAlHztGUyw
Dbho5UShAY3koTqDD6GUDoKVNAeflMyo89B5MgCY0h0NZlSuxD5LC8HyKeTgU5k/mXGpJJC8GcnQ
5lH1euMQiKYPXtRwtrZIPcrU0h5FKYnH0Xjzkv9Wgk3Hrg8Xs/EXu4AyB9jWPNuS5L7d9C1jzAe5
198v/cb2G7sROhBNnQUCtuAU+4516JM8LM6xhzEgrg5i16OFzBNOtnuvouK/HuYglmYTnJRd//y6
eJLTzHY/NIp0mdDlaO4NIacN2sr5iluklo+qopQ4i8cLrZM+aWM7bUhPM3uEdUBsBBiAi0KhFTRO
SVDAfH49SLSULjuF/lCJVEz0+jfGUIX8a2JNcsE2cpCnorrnIg+G2buT293Mj/7ri0f9pojEl4L0
ZG02glqjItfVUhHm5D/yIHbZ1hxbxZfxewr99aXqIVboUD93xPOx2CYLD+VMS4wQjiehUan63Zew
YYtBl9PuzVqzpvLF3g22TNKwJczoM2AoRugUW9UxzduYZMlRgDUNgk1jxlctt3oGeKQvSn+YURVh
w2npt0QhdHWALYA3/lANsMRoQpCUtaP4JfOPg/kHXh0EwqRPHDh6Yy5JBoXUocYlAwoNqBvh57fX
LvmZC9WyxPAaNgPYFKHFzxj/M7wulIGMrnk/KfWZZNhPwvvp7FgxORC30Po3pns9iPDbBip9WXLr
CpM0vOm0WEjVrHW11rkagMxBiIFiKn7LetT58cjTVqwBIszsVr46uKbFNp8x6Z9x2TREvI2KnuKd
ICSO5jX2BnApYo6ZNa3MGJ0SNx3fvlMvPuCwv7hZp8dS3Q4vZpOOrb66jFhw3x82Zm/mOJflliSO
5JY3wQjqZcRt/a1f8Dw4eTeBJF3PnJHIbCMXYPZNwmqhjHISd4qcOh8RXN+uXaFncD1l1+MjN/V1
O6hJxsvd3O7pV8MCCqxro442WHo+fo7jzO7rH9mCeGtClNO48MoSJ43h/DOAqrWS+KNNGYHe4Rmj
gm4NPsrDm4Ty2U4KOvJ85H6jQq61o3DH4GDPhAuqxT6dwDjHR52KVtz2RroD9EH9d77sfJxWrn0a
83g/MQU314NzmfNWGmk+6z/+Pf/B5hn07kkGlj6D9wSHjn5hy64ocwpqSXT7DF4Hs5/72cwSl5sC
f7aynXATMUiZ+NeAOakXIezpmr027MOvXCI1z4UvspvUOxLMRsEyVwLpYm+RTPZC2mJi0gotckIJ
dvHVhniTy3tS8XuPHUHkt9rlEnqS6fDYv02jxMlqo4ox+P4pQ6CVexoV24wRfVqdzxYMLGKDQfSi
AXA07oDlOYbyPx0RCPF2VXfv+rVhPDmZrUaDq66ZYUOb4TIzLzIqDYy22pobXhUhX4T44z7tsdrp
Ie/t5myo6HRelOk8sHE0+me4WlqF+BlyCWYtLP9k8Hkg51ieeGdz9UVYkqbzE/unTBfhpIK62YfG
iDsBXEKQ/LYGJh29jxyuflN0lglzmum9QidR2EAmo+/fXEeY/WZW59FqwUVqh35kqgEWYCVWe8E2
ntCdLnCa587XjgP2w3XaErmufeQZj4CLG3ajXY/9Nsij2Edo5xITRG5PTbP0gNL4Bx7/etG8TLO7
chH4TRL6LM4y3up5pwxX0Wk+X6Ukq8aquIzfK3Bo3vInPeg1RS24eYRqD+r8ir+bNk/Uhx46yGKC
KLRkLYOAYEV8PLl6YOhq+hszmEzL7Y8hv0ZiMIOCIEEp/iT1B7pfG9N1dmjCTWPYtHY+HXK/c2ac
4dmL0hMk/uWpozUgP63cKLb649UAk7iCCDpY/ovFIEHBnzG4Npjujh1ROX/cnOWfTfUTGtlWipk7
1Kqy50zMkQ59FTt+4vStaQaGlSeW4kn30SQxS33IRDF6pk3BUBiFvQf7UypzSabRaKVsHNGcSOFR
+4whHiOncGSxRONYeE3fkCXNbEWxi55dFEyWfbCOxEyk/FEvbk33OpLAJTIra0STY4iCobGjBQQt
mbFGhMehQhl/l5d+Ra9fnqxIBMXQhP5T+bWy9vUC/0mYQjCZmueVWpSy0/85yVKOEeJE2JuHzPu+
lBsuaQiEShs5mnf5+WZL42U4R13twLAP8ZOHFuUjCu1STsRnf51e7/mLJ+vqX1D3JIUJC46vrn5m
5CeeourXVW2fy9rkbV4OHwi94xLtLCL/T56b3uUSqsyB2xbdNPrrXxg3FyeLpBvGPoZ8mi8WD5hL
dK9AQ3yC5Q1nysSWWRI0gvN4P8nCjyylWYo4LItuTSjLD8zpI2X7xEwSlL5ZgWDhzkR70MPfi0zJ
/5GQi1F2tCAMNtAaORdvDHYstpgCEDJ30ZUJvoT5+yROUch9SnAczootT07PUVjeqJCp5mFMH9wQ
7Ltjw+KuUmEQu3vWb2qItwROp8tNc3SWcbRRG67mJ5m/5ZdKOovelYmZ1qI+fEm2E7J2N78QneCA
s/myKLFxxTPHGaTPyGl5YKiizRnnxVNWjfdVZhArnU/fJMgQLaeUeCeYu3ylcnO4hFGddxyt1fG1
2Mj0Zr6dNUMgX/2o/ImAWFfDNkBsFqSqdGk1xD35myakoHgQHVP8bE/ouf5JQ3HTfmD4req4Kbrd
0A+eor7epbQUK8VoNRkQ+vLbpRiYBKE+WRgFVhpI/VOvl8PFYgVWS2q5fylACd0+ewSLnUdE5x5J
+2JgitvTctBQ4VdevZqG80DweJ0v8TcWWVQ/UvmcKZHmH9xnQUGQ+OoGDnBPg7nFjSBYSwkM0UnI
MBxX6gki0mSkr+XeL81BVLpgjjqeauYQIF2qFWWNjFKVROTkgAVF4b5Btb+/LxzKrsuCvWByi+7s
taFU+eVTHC4lciMas8dfrtzjMxpUCwb5DvQpW9tTnHvtacqMnPJSFxxF07oWzYYj0Tgv8bX6tpzM
2SBVeNujgkBxN8fOH2SUZx6QeE3DaAvIohlzkRgU96lNgLv6Ci9LzphSBrYPDBqggX3IDP2sFySR
8V+WV1FKdXqAML9CUpFrECcySqiNN79NAiOCo1KK/wRktIXeAazYyHXF1bnfuYarbOpTwOx1isUH
T+xn9VZ5vDrK6hh6L3J1pbB5Hdjut/UQ9aD5A8vFooVP9O1/qSSDJo9BE8k2H266/y55aS1264wa
1lqhXH6cZ31aX+NXPC33ZdGn0fD5mcx6l6wPy3l1ds8Wj16ExKmLcqrymvJEtIJmxMvaeEbufdqy
IzF2AMgNPg61XT13wO2R6vBP0cUTLjJiHPuLRCNNDaX4MiIa97zxMDG3pXu6W3utLjK9uj47KZXv
wueMofaPIEWqnBrrN1XIUQw+dYmZTXSCmfCZNGpfVdjgir2ix32NWV0m2i0mr7/M9ySOa6cjfhvG
dMSoA1GxPVsAsKdmdSaYHo3tDq7dCA1FLPEhPg9MGbsc/z51jJcZg85GFURLoCC8eIXHZnpmZZgR
5oFFvKHYgJ6ntgpY3THxXu2Q2CKak0McZY5fRExXPVMJbxlG+kdfruQ4MtfpOmYndbOGfZr2Jyu4
6TiDeLZAyGFGZBMxA6u5LUicNL4QC3h952XNiVq1JACdWHJDeUiRqo349lKiqnwFDN3djFC/yY71
Srg8jNZGqJUJWYS5uXmxXj592dcmkrreqHd+v3WKg84nL96owGTf8h7Z5hH4+3RYVFnnaSjntWVv
slzuSTe4nKqLG/P6lPjdLlBC3xkjKw1OOQ+t1Bh3/kIDffxjhwVbLgLOvZEZ/Me9CzM76m765yqS
mVKLOAIGA9VSCfs9um2EuzXFaboctIGL0RGEq50ud5vsgKp7qYEwwljZ3YFXTWGiNrzvnn4EiBHf
IlN0rg2HlbUTzcjAwLc6Utz1fvR506bfEEGi1qClSi3igRkvhNzMvB+aTYJ2eoEU8rfX3pTZIItV
xoxXWkw+L24PC3kAT2Lw/6SZ/Y3Y9T6DulsvNqyGXibXJXfw3n6m+W2NrBmMP89yHKDI/ihlQTO6
fv3N8VSR/7weIpgMrm6+Zmar+84BanY+4tA1HlFdltLVdAUDH+RFfeQ5N5zQBLWgZh+FEw0S92TB
TLH7/aZsAtBpQgTm0YONXU6Lm9mBDGlwndS78fa5D4dXp1pvkNVZmy6RZen5IprKnIQ5CHTeOT8f
dO8btKESsYPPnOWFGRiR8ywC2b1JDUgZc8ZzG/eK/j/Z21pOrhbHyOSt29zdCUhqXNfaPCHaX2SO
BikPmBEfJPLhMkakgmvn56omyjnSr0KL/b4vw7dlpv3CC/7GRWETRvUvKU8eeYWNO8MjsyoOffOG
E7cKoR8BKOijubEQ77zhpT3nTT7UmV8I+NP9AUBI71zu5DHhUcNqFPvM8l9OiaXZnYJChnhNFuzh
9TKUZX9yvJB6QGVTYhqvYCSMPR/4HBv6X4yULFxnRXwu/QbPhdUUSabpU2LDJcpdWMOxo+1GYZOj
d2TfvD0aB2Ayc+8nNkuYBXgwBSY8HqKYnJQQ9d4xlCVKv1OuYpeIKHLB0gf/HBofARXeqxr3eEpZ
RPpK3ooRNESVgZYMyvL6GVl/p+3H7rfKjhdLvOvYE8bVmjXBsVUozhpyBTbfKrVz6GZAlU9rtho3
mZR1tC52L+tETwghGKRr3qVubkinWeJxLATSFooSnVgjQEk1XbzMrSxI5anhr0Mzd9jpIVd/jJ5E
AIM4hDfQWnX3ZDweBohJw1WdfL0QKItC/a4CwGBxFQF4hLgj+TPnHnVh5yHne3u8QtAWLY+gyOaS
lEF5GhVoDMxvJYvmA/mjRfg/gXzZyVs2vZEnKAJ8MPKT4+8apOXbYrxgbhu5JrxwRFmWqYVa61T9
UcUHNB81bVFFulN+7BSzHhJUdkRFQUCNj1YNhpBGKkXM/V7+hnUQ0z5af/RSrlFBmHPa2gnvVZtx
BoqEYEczT/XMY7wZlxJ4KIdHQibOq3xxtZ6aECGLO5nIgzgAu+cHP1AHeovjUj8WBh5EvC1f0Fg6
wHQpF+F43ssxLCLY21v8OKVK6ZGWEjsvQN0at0S7jec5TOoZCUa75/kpXQZGv/GGAxkthqtBT0dl
FUeDMxRpHMch2LCVem87x8cs5OH2rQPxbDJeGO4mC3vaS0sb5ZSkLGouae9LxpXxBAm+RxVHnLpR
c+A1YJm/8lbXOhnSI2YUyBy0FgEoh89hSixWraQe3JGlbrhIJ0OY3h1O7+UnYzTuydnCYt8ahOUe
RAkYoFt6koxG6KWU0T4trYBN5i507OmH14ehKS9sUJvUWd42gfqd4GU73vsEOIQHPNhnbi7toV7X
/CerSYygzzIk9YG2R6SMm3+RR+EBZRqE0MBO+tZXZI1r8hsFWZfADZK86tPqxJF2VMJ2aNoSjJmM
MuejI8Kl1KZsz3byJQvs6YHHFCLm+bIllSU75naZG8onOpDiVZWpM8nK2kl+INUuiW/uxXivC6NG
r1FeZSA6v4oE8a3TYln5N+WpvD7M9DmrRb1AvNUYawk4OQOkAKqswY1TxlJTEpG3vnrHHlgZf6bV
gguoSGqV11OCZg1M7T9D2DkxpNIAdcLccV/nwF5U0zKAJXMBNO4+VSwVhTwVN8xjHiQQLF1UJZYb
yv3Bi6dQd9nC/9ERUtAfWStjUbXmQy7P7aNJicPd18QyMm80nO2kper0y7UtVzJIiHMPmAN0gUjy
DD3RsTnL7RrrBe8nikAw98rWaFSsbebTctxQjZjigaz904UuhksRf+PJ69t63a6s9/jZZnmRMADW
EYt06C1ehs3O6/y8T+zfzRyy7OPzZRQNnbGgLVjRUIKuPUKwfq4Mzi8IbiJGkybFY4taqi/55MC3
/tFQAUv+Iy+GS8v24Ndc/0YP9SuPFu6wEK4aeXFm2gTYT0oF/Z9GDFsrH05MQSXfaLOsJKXfgtQQ
IGO37jWphkxewDxtPJ/3VPB87DRv+Z/XCwILBbqHNTRzr4Kt3/y+j5uWqkU2X3iXvhZ77Mk4Mruo
gTX1hTo+SBdcNxi17tTdW/hbNDUvxJ6tX2BjpEMekn4vKPxO3UudCM9r3ozcUu2VRLlNdUqznXE4
SgYLMhQhw8Rh3/wNP+1d/I4sH2tuOnDbtg8wqLfIf4eVOkGkpY3UVfj09A6bM7lVGeXFZR3ezHau
9o0N0dcrU3oe6LKszOI/la7V/FxeOaJG9+7+S0m3nwUGFvh+APmlp55Od+n9mEPQPG8B05/2eZiL
NX+dCfyuFecoM+HE4Sj7vQhUNzfHQ7ivcZSlLE38FL2HiT7pY44lccYn2op6h8KZN3iERWp3GKOg
MIVNReBoQZKZyEfGsV5TyJkf7EkxyHRGaaSPh9NQ3XTonxsmOpVXZspoMLSgYIorAYg+BDDRDAM/
SBOaLIu5XxXWGEiCPmVmlsf2Icd3wEyhYNMdaciOXLtooP+8u97L7fr419ruBUnuDYm81L/qzeFx
Dug8O9JXMLI6vfykm/LFjDRVDF2TahsR2KYetPwzzwOpNlf0WTzfa9jdUql9/S+vp7bfSk2EGC21
W79tECxpanvQrOT/Uu/vZ+kEETNkjvnnlxJ9IVcb61V5croZoQe+iRzzhxNFFHwuxvRpg0/4OeNV
TnQ0rIYRIebutEFiTidActG5xoamK3SMThMt4fOOqPDy75lMibns0Elk00tYYrhd/okQwgr7GgkN
gNJNytED6nGnsocBk/LN5STM68BSMg3datGystwAX+LZah98vCSk/QFmXlAkKtpNp51dR4jS7HcN
TBgckHByiW1R1wgs7aHdIOPRkqBdtn8UPcJ5pNk55uiizA778HNCBiNM360nVN43rpSy475w8KPz
EJUpFIE+B1qk6oz7k/MpFqfMX2xXLG1s5k6h4RYvD1QFA+E8WDhu9WvtCU0iz12VISZKpxlH0kMo
9u/Ra6UaxG1kBzPNlYNqhlkFg5Hy2iL9r9NmRnEg57GePvJwxURZ9A7vhaM0WieauBQV27xCGgZo
jlr9kgcHT8hGF7a0cHYSzcHnWnDrzqsjgm2Qr7josRm4f1AmeAAHI3O1scdBK21ZER9elFZOy1UA
upwiXUV7n1+hr/pa6rfL0fyBmsF6vFjv/qyfYtsPjX7wd117F/AfJRoE1lm7264hoIzJMEVSQfKc
FjptosN9xBk2qRi7Kua+ccQyyre4HbTS0XvIvpbAn7rkomZd7+yXrMYvQuuWwuq7i1iVX9vTuGgq
KuJiEu1cG7vfujzMCobJ7RGjbPI6ZouPdsl7y5pKu4NwcC5gI7tqeufPFlJZ580+gjoAWBGQ2G6w
0v2Z4SipKpRcXb5K/hlbMeW/R/ViXKRq2h5//qTYOZ1WXwNIJj+St5rGFBsrj94EPycsQKyuZW8N
CHQ051B5qVho7+HFgR35Gv0mqKG1ZypUNZJx6PDTpzqSRFA3zzUGVuiHXk5QGnwW7Ead9jkMulAr
sBOiKdPE/QRO9iukQ2P2UrtIN2p3B4B2qJxjKqreMCH1MRFMJH2eSJtNbKrn35VmkiTnIctPEq8F
XNKfu/SlJ+v3CS0yLh2g9Ckwuyy4cWrdBN0J5WzOvKv+HROFm06dXunjPWEMgF5ljb2KGck3qh4o
qpeyXNF1jwqcSQCm7eMawfwfjb0wTzRu70ljItKHJkKinDnOYlQ8IO7/L7stF3RU4GnwaqDfFl+I
nPeB9FbD+rRI41m3QQbv3zAeuQYItgHkA/+Lm0l11+rMTUkLpvmYAwHwx9I12kIr6pSdIDQ2Xqgh
FA2mn8EH0rBnkAeVufJOvjJkSn0DnnqpCAgLLnUYX0j29oeE745zqmpL0gPH9L4fo4dXkikL+yZn
KVM16gouww/GWWWMPgldGzzDdEPISaeTGMCvjC55RYmaStzHujj92Pm0jlSijRFU6OYIfUq+nkkf
nMKxesNmODR7Vw0DHE8co2EAiquWJ388NtgEsrHsa1A81v8LvtGqmC2A6i+08aLE517SWdwA+gvi
meh6NuN5OJLaR/xcpo30MN35mc0xJr/VOiTzh8ovoWzhn3uWrgzI0XOhSiu+AHWyN8mElS+q7Cre
czrpFbSkqV0pVwJMXA+CkpN5DkuHMtyVkmY92w4XbVl+x4liCBsblk1180yn5gmeiBNCEjyfCkKG
GnZ1XmKuYA9n8VZGdSGuNVVSVtjk1ar5CQbpJzYR0L6W0uo4W91XlkafrgT9+Rt3dt1y0kBM3eQB
myYxxD28MV3zTSCGliDsKd0DThNMryRj2KRf6FMq+0ftJSxGgOoCAnma61NnAXInFXvzyrE/9lOT
kG+j4L07pdZUOup2tSTZsQAlx6M4sc6rJtK7GHyYGidhUWJWzUxYEUFec1KgLHxBL6/ZEUV28kCI
/mgYPmnwbYw+5EHTMGMtUS3evUqxpjZ/bMmzsc2YGR4zvm1PtcYzY9ea/hXON8hHdYxq1SND0eGI
7g7sijAfGQfFW/WwMcOFItIh/QKaP8gDLBxgIBrZbgJQMihQSCjcT5msf8GfEtCZl5G3en0FQNie
nmONtG5fM4EuokkOEhWdvPwndOcrRJ07HLEWSbSqZtfz805vm4vvHTByPVCn4jem13nSdyOyDDX7
gfK3AC8NKDmCEaWJqR7TKAI+rx26HaxugnvjGzwiY0GYhzKV4ozpeJj3AAaQbA8iljaNeXOb+AI9
vRLZHUgoF51AKxRKPgLpEoId9b8tMqKOOTNn1yP3lluyE8ki/eyT/0AXGO9iFa1uPPtvHHRv8i8M
TeKJVUEvCWru10xAEZxh+lkk7gFKWGdCxGBFNI4MXFEXTgZul4SdsxxVdFkrizrULWc3LBsmOWrl
tzZRMEFcccJGPFYiZYqcY+cxRcaIbGNzp10mzHvxGAdnM4ZLMqsaGo6MgpFPdA6YsX5G/DgUhh3S
JDjDFQyLRqSwqKjAncZYx+jcPebXonSENmy/JReZY9eNsIRIVJhujbsyFTmT5HtMQMsEvP/cKTVe
cj6sIgr/ljdL7DytDM+Z2J8pXrBRPoWKKtcqt+TcUJtMBx9XYKELbXr5/yJRvdZRq2KKjG4Fih6P
JIBPeNQd3NHYaXE/yY02CYtb4fuh199t/fg4kXRlP0Fq6cP67cl0PuADU2OFEy4uCpWru/57KMrV
4acJM3lGSzRdrrAK34XXwVzATEmYb0z27pgtodnlv6Cj3qPE0GEYgMWF5tCdNMs+qlBc8xa+OZgo
6v+DryvdVGq3uWmZdKdDOPAzUMhvghAX/FgWNei3bshCe99ZMR0lh5Di7EK4Ngo0rvO9ZMNAdo8F
8vfqd0Cm8ZC9DbiFO/mV0pZzM2B/I/8mkkBfwvhzwZ5TI30oZIrMJ7OROy+udFjNDgt1oiVZXBQe
bKyNuhSpLhvNbBr4YFttuEv86UIS1BGorIZ6G7Dvr06v+Q1Q+2zUzi554/gTpNivBWRrFPwxhsIy
zjEFWuHlN0b4Xlm5pdTMg7Ha8E1otgc2F6Jus1PAC1EQ5HTvjFDwMyaVzoKEr8KrvDngmfg96+rX
I7oOOGAizsivdXAN80vhxmlmYORSiTuWZHtS22Dh/MTyO+yiBeqGmn42TxP/ZEf8iR9jmmn8zs8v
HO8Il7xYpFU8Qgc/I0s3YupiFkaAtGi4kyaN+w527+A7CtcRPKTdKGcDe2g0adjDPJ1IGMWt9ehN
mdzba6NGMn/JbFXqNzRerKW3toHEYh49eQyI7hjecJYIL/r2WrEbRWkjGd/zMSZQkGAjSR/klhKH
4AmNhVh4q6OXUgZAOnK1tbWBnMKwDWbD+JehICkhnNoAOzHB4de9c7t6cD1gAW+1KjHKOP09RIID
vuPD0kLsFeIMs/NACHnbneHIGCPCRfVwffBTIyPcnZV+7xzRh8w//im+nISjscODKo/UOVCu+Ial
Zz3ZX1rBBf7hkDq/nyos0fxHBEUOcT4O32Ox27uXY2r+SrZxbfLtM8AJzHliayiG5bv/doHjjJYm
VsDL5nbDw/OGPqrrIquJotV23DasL0JwcUt5+bil41JW41FYH9gRA1sJwG21dIMkNjqZk/Wtt2pg
OX6f32bDWzDaZrzE1RNI3k0XdTRPM6cBfsxRpOivcnFuTt0XU7FoI/M98ZdntRsJ0mMldssICHqa
BVRFN7D+/qZKXRPZlffzjPqejCY48g2WBD1bRewg6UCmWeBOXyX/BexHZ8mSWGsengDcjlvYnSWa
aOz5tj/8QbQAzCSHeurt8PQ/muqOYLZVElz0s4dLWrnhRXnjDWlbvlvYtWRHpAtvQxBEMd3spC3R
dYnyhSjSh1eAkn7GeBXnYguIvHNWTasBlfbkVFQb5cDklRXACvjomwgvMqzCU3HSQgPvld+P21JC
3cbHwfeylIRJenDvhnYJlvHgNr4CSC7kk8jKIOTEpZ9HsMeCVN9sL3vADegEuBMuk1MwIMZH50sD
xdgNBdTIXhR/642EeL05bG/XWrhls1flDWTBntzqHixxDf4RdvEu/GJ3bKge87N7hZRFQrH/QYCF
zCYGwfyBd29ypCsnv8kpXPQMcyQPscb2/l2SGAF6Gx8W5RGb7xRlxYNMOEEnf4X8oon0Y6YOS6Vh
nKNm/B7C/wvBTANEglhHakV8Mx7Bg9pGpZE1doUyZM4X0JR6gpqdQf2TRCOl5UER7coQde+QT8Ae
/FzVbMFCJVMlGrhW48rSkdbYBgqRHXMVen494e63HAKUv7VdZ5//Xq3+L97qM/R/onxcJ/OaRqqX
BPjPzc6MZrR/f47AfTKsDctZ6OVK2f/ggk4DBh6/ZDvIuznK56VyBkVM+Grx7WZAoFrqe7Bwo2Rj
FrktIcHZk2UD5FIcs2XrsHT0LHmE02FAhOvoS2tcWDKpVz34ojqGjhFJx8ZXO5B50O2mkqZqi0A2
QjT7Mp3ECBDOaqqHQTxJIfTNOqTWKDAFeS0e6VTxdECQVc/otkJIfpDfDloYJjMn2ljFjsZdeGRN
Nu1HHuHYkMbEoRN397nJ35ogWplfsU7zNpITG8wlgT6pRrBglHT1+lIkc65+Om9aRvqleqs0K/pG
XBMaAHxV8RQy7hYQc4+yaTBsTpvcN+dxNosa1VWFEqr5to+G0cSVKoaCb2+u3206OARtNHNbXVh/
Hp+bBOtDNVxp2iXJPnCje5HKk89ugsE26IvRCpXCohVaZ4z8WXmRB0+pdNf/SmfTZTbOmFkJkREo
vpjyFuMTbpHdYXUprQ7OK1hUevoOZ1i+rwe9G4ZYcsK/XGYN9FsOKR0vQB8P23M3N10XJD1Us8kL
JXS3DmeCDcBfoX+Y0cmLELjMvMKakk9BtPcHFieH5u0gSRpnOfY06iQQPv2OIK5H2lBNGbuf4Xzs
jvBbprxWuj0ie/3WUV7ofj7/zp3RhVkvCnKGSwU/GmTiFVp8duAK1oZjLL4GThdCIznggi7jxY63
XqkfJ3FKulejJcpztWIRQlybcJfvpVWNo1s/M2W/wKeT6m0lQjUNVR7Cimo5j0a42o0SUfz0Wo/T
G7OUp97cS9hf5b3wMGGYVhddyntFQ/YhIlpkYuz1NJdLVwbQNsYtxH4ovqDVYecGalPkpAwlQCAe
7P6O8k+LWXGtEH2/zY2A0CNPy7SsU4RJLGPWRcSjYefO81BIS9RzdQ4xAunRNaC8VKh0IBJr/hDG
uiV4gC85g9QrkGkZWeacMF8UZvcOTI8jDlvnCAtz4wfE7AjMh+A68R5JaFJSvdxgG4BJkdlVKJxz
p9FH/Bm636C1LYBVp92NeDGz+5S+mQYCXmQ/6yFBMjgWL0RZ0o5loQOE35NPUoW1jyGVQ6ETGRzJ
yzCLtLQO3nm3Ao0taiq9sQc2msMuO3X621pntNxiSeJDyNfHzvuFdfBwBUWKa856RSSxVGKy7r6b
mE5ES1l/JKv54RNlmHCn8cFmGE4SiLxOtxNVheYLrNK6RxEKWL7yc9EVHILa0iFEPmG7BMq6MxZ9
v6OK0DJx94oPugFByIzTPnNnjTv35133ekFX9eMqafPSRJJR4bgolOlQEDtilhhdHKDfajS58DZ/
K/duA8awZUNfx/1KhTuYnB2V/yJpBxTNg1BwYDKHykr7pfgYcYgrVlSq/bj6jN87XhSHGWg0GEJG
yh/SrTMKDDWwwbRZc3uBYQ2n+61KMTlC56a4qXha34gGagU5yQtgfF2Z6NRud6rSWSUI5+GXOis4
sEMsQ2A+V/OldkH1/K3GLX27JWhK0My+yy/CEmJkb2eLrlil9F2hi1TaM+nidfhCv1mFOgsiQPXx
gwY/4p2/rWrHJiF7MMtqgoSoHsqhyn6MKUEbp/bed/P1xBKjPwjIlvEUPJLjVcz0lK2Trgv8Igjf
jusjQIg0Svunu7D86kgWWVZdL7TsThIPx8qCBss/qZpEhWqpEtUKg0p7pqJ6czBFnxgtOPP8tXL7
GsOCIHo1Z3pn69zUMx0+EQHDerLdnwmQvlxWr+YiaQiQeOoypnMG0tODExmfwoo3kwpo6sIzK2Za
VBzGyw/JD+7hc2ZwOpl8HKVXMXadLkxLBy7Y34aTonBMxT4ELmOJl6Pa1TNiLzA9vU6UbD8fwKmg
6sz25AWixHw6/smQJ33U4TR2ZDPmjXD4SLYW74btXydEJHi5cft9AQvgYMwAYE2BEFZ4Fnhxh8YN
vjhZhph/cKKG94aL7bVMq73GhXD9HULPHxEhxmj2Nl3M4iEUt54VFjYCN3Fy/8E1dVehUd6PBx9V
8kONu/FPkwVtrhNhhANSJlWTRbG2E3JxTfkFM9xvhK1DwDJUqDO66w7oQ+7kVj1ruJP/wiMPr8xH
HJQ9qLOwSvaaopAsn1WFsvnTGSfAPwobqZdjXKyNpQHMMYAsWi4hLsGzRb2SiZteswyR54MX9A5Q
L0woowNMTMHbf3AP6fxMP3dWMUrFBEGJ8nX1AMz4KkRWdo9EmbA7dAmHy+WNq+HWX7wF5nQU/qaf
QzUKfHP9ejc+F+ZyYpPkrDkRSJWyCNvTwVlVrwn3Wn5Var+vgtIryXYGoMqAK5HZG1uJ/wJUmDX5
N6ShTH8gL8+HBK3jMusUrKCUvvk/Mejjt9X4s00NFQKL2/A9DrxDNxuCCmdR5TlemHI3vK5dFldd
wInefPr77FIaFh2nDESRQgUl2zpu8ltl6WZlkJkRgdoFn0gtTh0ajz5Of5UJGd51Z6NZT2ov0suF
+HHrrda4YeY2xRS1E951zMUgGL7V6L2O3t2dM3/RnhZzm9IgiBehB76pZyBoSJRD1IMwufkDRUQS
bgMWZ9SjTKZuWfJYXM0xxLC7FEqhfLIuTaDrDjUjmyyda5fq7s8sxwHRwGNFxj+N5RiDwPdcD6GF
uPnG9pIN53PV+6k5q0yVEpTdj77OJLkEZ7rJ/35T6EYigt1s3UNdchwwHxSiy2qLoqWyjWzsPDZI
RRpzxfu5SexSH84yrS++3CDnL66PBUr2VyO0HtCX+IvDWc3HDFdFBt0+OFx7Z00I0mzuiLsVLOyB
sUTFGXFeds2EAVwjOcXO8Z8OUdLObDopPI+oBYvfcICMWivPXGU1YgGHDVq3CZD7Dqouu112W8Rl
QtK205OmBMiATCfRmy3FsR9wQ3WaJIBOklDFxZs4t3iNQcbF0JoeeCePPb/n4blbWEugrJK7F1Zb
3hnkZg+Ew63aFtvLWKtn9wpScCsqAhb6+noEHl3WPrVVSYisAcDerDVQ02UTMPohk6L4MqE0SwC5
GLxN0ph7Es1B9RltbKgPnsIoe63cmm8rbGzAWPpNLV286uASvXH8e5SXx0CV3QHiTLT08tkOGP+i
Bwp8P1eNYQEr7DGdBlbbbvCGSjwhdhQ/tFKkkE3ODUbbtvW73K0anoj/0/3iDAxgKOLjb85xLKaS
NxH3BcnHA7vLJ040ewSGyRybCSJdUAZy0brnw+rW4gmTqGPLr0nNal4DT7HNZq4ygCoEdeQ7smAA
RO0fwRArnqiuA+K0woxdL4798fG63Zc3BfOKhIBNy1ecqLLiVvqp6bWB7BNNjdURPMjYKZNKek7V
hAY61VH6+b7Jn6I/+lhAELMfcY7vD4Tuv+2Px1YvqdoXK3RUDAk+dTHOnDNoyYdkUt+aS04zFtxL
pDLAd1YZvzZh4R/R8f5NFQjXSdrliPcF/Vjbk0f5x8njUnb2T3O6FkpAp8oHREMXyBUYZwgUD4T/
G8NbuT6OzHIHm8MtFI8slxJNmdjWiRXIrU+joeP+Uy0N6VzHyOrBWvtNNgw41eFtYeT4crDPvc5q
d0dyO2HQC1+cqaOD9se5G9DqmXWEEiZDmdrM7ssJ6GwGRHm8oItkFQBNEUNOTugPV1+Wz+sBoWRz
hfymPRM4frKpx8fPFx1aO1NQsrgVTEt3yhp6mjJpdQIzcQlVfVc8xz5HuaTX1UhJFHihzNxwhj67
0X4a05T2I1ALYL3ok3pym5hnlK/KYYSeBeB9dEC7LRN2TwFnZhYf1TQrqn6rnBRfuxhU0Qq1NQFu
9dlFmGctXI9UCJTcYrYa7i1/3vgYVBVbScnfuUxS4xpofXtEWCHYoN562xLT9sx6qpIwIAprWqB9
Z19ik9dEXR5sWP1BbSSU8oxJef05KjEgk6YQPycEQYTNOtEUixzGfOEllBOmBqIdEy6vJsc2KHXF
olIiQ5+YMkEvi2w/SHHJ5wBH6QnS57uP9qjBkPPap0FgfQCJC5YJ78PLW5yiqpy5Ggr8N7dmhmlg
UMpFDqsgmIeWTVZHNv/B9cisz1zQVTF7eZZ93QI9TXwZrYbgeaFxgFooU4mY4XnDArPohcTtDTub
89SThsDYWp9X/c/RBmMFCgvyCFSEifyopWSnRqSxoTIESwUOWnrkFQ5A2+sR7QtylJlF8fCDohU4
QPEQEj3RiDkHFTIWyAkw5+XHlQUBebYthZL4QXNVfuIq6db06gGCoV4XIPXtGtWll0YCgd1ZtWL7
oR52ieSo4tIZR52k0WcNtLJgv/hp8CWLFyisy7ri0/Qr3aWPIsc2jyvI6LrlLTOqjHe0Y2fe1DhQ
QngtfTbKBqwOZ8n46TyQfvaJ79XG1Q8W34T26FcayRI4PNgWnhqWfPtSf8oLEHtZHm4vAvah1cMi
Kit3ouElbli97ViqBktEBbzkXu0318hPpUL2ojSlpDEdOPEoDcSVFtN3mshvtLVJKcDZ8rbjozgM
8bfPuBnZ28n0HgYjO/uFAXbMxxhXjxXOOXKEfWsNPVz6glLNqF1V6CZCUX1twUuVBDLE//sXt56Q
+n8Wcd/MCkqC0e8/97wrA4wXNJYlzsmJcjJduXo7LrlJl9WIGMzcwLdcU615aU/AQYuhozDOWsts
PVyDIEMni9rX4e2asURWKlcsCOEZUuxqnUIdwaHsm8jOdpiKDtPuZIFuYxVlXQb/aYfEw5XK9urL
g4hVWGZemKZKbbdsb/lMXiV3YyLtsJV5JL+s0SPeTyOSlCCD5sSFmKO89fTyHALm2MacBjFuQuXY
H+eJrRnYYVj6m/qt6M7xOuwrD5IML1Drx8Tq6kxrN4JE2axG3kfEThRAinWmlQ/VXW5cKS7mk2dh
fidTepxIeeokakRL5A7KbvUtTWZBdQKQoesRb1BX9g+0qQ8sQR/9DyS0Llkh0ED43cJObUOt/+Oc
Sm7UT0yim+U61bMlQDBt4Wn3RwAnHKZZ3kCRlXCOVLANnuBT0kMhmcenMaV3ch3tW19nb9O+Z9xc
8KRp9J9SUS6+OyCpgglJThJimUL+j4QqXSwJueMNnbVeNMTmIeq9CWJh8GvW8H8HtJGEFW83+TFg
SRZ2fZTyzllyiiwHZ9wJih0aGcH3VXrdYVEutWFQAMHkH9Dpb00P+afTSfsz5DkTgaqpeyYYri1s
Dz3T7zjdSnzM1PIO9SM99mshbIsUePERTPNwOECAtFqCovdNSmz8QHk+clQX+Xsf6uaQ4I3cWLfj
t/1+VsevYKCEf0zCMcgLOGaCsghKaeCBfO1JP4caQ9Hye5EVnCWGOqpqhWX7OpQG8xQ8Cy5JQk2V
d0oOOHOoY+dBZGLwxcD0Yy/FWB3pir1b0vrQtriAYyatID1mM+h9so05QsmQWiQTi1/rWQvpW6Ps
Vm+HG1mrtEXol7LbK1bKrq+iZ0+ZHwFA5swsj0EK0pXQMxTKBaXZJ2LYRYN4pQEi2CL9y0M6V138
Ur96UM2rdJJFn4LPEr+6Ci+z5NmV1SRLoXtFxfIPRq9Mq1eUpEnR0FQf7k4eA3g9+YZQyDXOHMsQ
Yh9AfS4iPbvcsUtXu6gh737NhVh2p4R+mH9POnZGHeh+LRTY/Sks0H4qJ0Z6CvImwsNMxzlZPDII
SeIKAAp8a2BOqSV/rAURv+OC05X2lZhOcluklN3wp/526eIsUWle2J9CV0GU3VJ2ZC4a0MGEbOyO
0VRRwQjHPGrR8QNA2IHj4bWUbRnfHuzD7vv5sVk/ZGgvo3Rt2jkOEckM23KAyTpJy43kRS1UQX8W
nPQh2O10veWAQefQB3WXkco1JQ9dU8eh4aQx0MQlAhVCCWdUjxEk8+0d8jsdNbod4oqfCSIHNqcX
j5hzOZIh2a8VScLd1d3gRZQ4LjZdO0NZG3z9pYBWBhoVdngOH5D7Wd2ijqTtoeDTJCZjV6aYgOiW
UGLxwWXv+Sfe4KRvWl3UGZJQNSRZk9uvEAAOF4tkRvtBACH+IsiZzhAKYXrYglicl1xGq1VL1/GN
Wu1d5whHAwkWKsQz96qdx00DeH8AJDm2Yd16IW1VsjYUYx+meL19k2wr4I4Ybh3LNxftJRjOn7Nh
xNn2URUdlGS9ts26diQzDmWc/17nuUOquYHFfdiKSo/CvARolknD1Jnnls8rt38fbpdocpdIsePq
HydBcXsFx+rVJsKpTFNjkKtLd9k+CoT6D//d3ONNx96bePbG8oOOE4MLp6lTDvXMKZpOuG6yPXA9
h9yET2Fg7kWlWtS03bhzkkzXWcuqWJUb6C9fCHTA6sI8sTwugW8IStzDWQI/gpqoUTvJRStOb786
4pysx8Bo917oTetc94bCz1m6ZUR+6K/gTxAQ91iW2xPtte31sSSLZRtsQoTrq2Fp8G/MsOr6VH6Q
XVFgiS1JxsbQATngnjwDrbSkZHGv4nwUrJSC6m0ESZZgO9NSVganQ7lemRNtaF4Xx0Nla6gHMnLv
6cnOuoP9J7wBYkcgI4i2roT4fBZTu35zY1BKw32m4g0InKNPt8MLDDTENBGtKb0QiCFoQqYY3ehB
iUlGEdo4dogY4vs6DxERWaUGF9h/jjdHrBs1W3GJvpZvnssEvQ202B2xaFTqP76odm59eE/a3QV2
r7RztgwO3xTuygKNZTEeUDgk6nJQ4cXMGilaEGzpIvavVyRbuxP4FmSVWw8yAewXGs20JyFVc0Tu
osVbjtfyL59FtgCTdC2QOnUaGd81l+da0/LJ3GOvdX5r/zLYpqUk6lH+yjscMSh3DBrRQhLFkjUn
/edwxUe+p+8IjS1ZGOZGs5eDMvvgwtk+QdQDVxE/3cR2mnaW5bsm0ZTAh5XvJAjBUXFw+SPJWudD
Ty/j2iiFxGr+WEXovnCPb6vL18pf77Eq5EOX4Dn+qylrxbXmXARRVHP5D5dAWGZWRn7BrJKmW267
EcMHE8akDx9A7nzzh4M10AzCAG/m/M3SbNEZUq69iep0RNkE2e4iR3eJ4X7XsFnk1gtkJ53nVJTZ
e7Wp7F68nTPOfo+hwJ92c3i48K05Nv0Sq8DNczsl+GKYJRVzQHtxqd8/VsGDsGXdhr+ZiTd3fND7
2o9lvd1iGSZZptstlZm0RYEAY6+4ZNVwPu/kFw3ruLOiLp/HFneRxHLsabpLKy8KBAdEnWgrnvMo
+LYs+Sqrl1PzsWZ2Qe3R7aI/FjyD/4iRx++niN631W7i/sHb8YXC/KKM8J19eb7Wf+wL4UgkXWOz
R60p1pkvI/ThOdzyd9Wf4s/mdh47373Sy/MKzh+SCm6ZZ1xxCVpNuTeiZLLBOUBkc3xIgel53xXz
Jdb1b1Z/ufTwrjPO/wfvJxT7tFNhJHbeTyojxDZttrDvf9jWR6UAyo7f6d3J3kocCPuV7L1Ts2VD
OBJotOs+SICTJ//xE5A9B5rZ0AlSBCtqZPn8eNlXjMS+1+Vfn4PKD6zzD9d8AsWLSgVKta8Kxtj0
UxZrbmXsuteKgHvW7+dq7ptcsW5v73XbYCjKOkMrVMrEhxccsnlXh9JDBK054uF/jgx8sp1Q3G+R
W88OjUhF5Ntj/mJsNqDDxLeTJJfyryQ5oU5qQGqzkPmWwv8NCfIQJJtaXgbWd/GyJ14F4r1SOgxw
xDUZHc7BcRpU/hD1zTPx6PZPvqiTmY4x0eteDh0bXYWaPLZ9QOe0aCUFmR9Ea1orEkJnulmX4wVj
g2cbEn+LRKpFWrVJ65F1rOInelbJNp6KALGVA+LCxAcJWpIHI6QtIPuS4CzLDiXHRFOuCVIM9lGu
iQGbWNuDlm16d7N4z6ifBlTaSc4OD6SZRaZjtwzw0s5y0evoRYYztapSxkNM/mGkYupDAlvPkKPx
NAkadml5uRZJkra4s9E2RzPFBzk1wfudi+Ghx8Cot8wE9t9uNKlkIVy4MZh0Gh/SptLR9SHVI5rP
AMzhzAZF3JN7IJUXd2BOseDwxLibTs/sBd3oqQ80GlkIWfURbFxQuMHr7GY+Wit4nMUIiIwbnxiL
r+Lm3LfGE2IJOjCD/y3Pp51ajOi6Ol0yDjlf+Az6IKQhD74FpRBhiVneCp3UtTKWntCp3r+AX70a
/Kr5Y0Z+FJehW3IsAbxZCOlEF6PQVKQXFyNmG95athybl97OHh3EqRzDOm7Id3A3/vNaIS1x46qe
0YPV0Kp8nIB3LIF50iKGdXXFQ0YrWEEjocylRWsjsZgPcTT4WW5jvvQnxHaX80ZkfY0aBEFA2CU9
J5ukx5oTVmerlHyfkQ6Hn/KWZ7FD3Ae8J4c+QXoJLAf6RlFEjBf7vD7cxcBcnoDmuDhh7DR+7/A6
HmglI+ESOK4jhDwGPgOk4R5/glHpoVImlurESfP+qEQ3S59yG313CuaVabwbbOKw3eBTHfeS9R4X
RD/r4UEDspjispTW6MI8s62siYy9fk3hOQlDQ9jRshpSrnnPeSuIzNA67IAA3Vh8VUFKQX9ILkNg
HXvck7a5JSWYoUuSUVoQdH6GnypnyR5+mkupnhaJpbbEqZTTvAm/LQF87dmB4CV4LWH2HmoQBACo
YonYbMH11vYsvReD9P7V/GDNTKtg/qqqDQyMIuwCPzxcLxCf1dneiotMbz/pXCfTfu72OmMrjJ+U
P5Gew3W/m1MTQN22mls1oablTYY9ZYiD9tyenlw5u5u417nms5vK8AeK6M8EukjzvG/VrnAskml9
L4urOZNbeXhqkNJ5i3lmGSvy87LHBsZ6Kp6TMJ+3Q8/qu5P5EE/o2HPtjWBcTtuayV5h2PsuL/pl
EEmrQzvSvoe+RYBDkv113O0NFDUZtjd8qd2GCwloz7CyoZlAmfQhsZHNFZoERLx3GGniFdDI12RI
MrUqBFHzfNyca8Nhfl156TX49YOAffTWiGDreZRrDltvWqJ2Z9mBGnWxhu59LjFgvTQ1FOTQPat1
lIB6JOWloTFXBrVhbFIg4lYpWFgUAL4VC6Piz2IOkl+1YE1kbHUmuDjkMCYk3UBq3cU9hT5Bsp7/
XUioSFRMMUUVtSVEdIV4fuLJhpTC4WxXKvk5gU0IZqpmT3o4bevvnzQyLm615s6qI0tbY5Nh05/n
uAdo6E9liPQpzgv1uELbDWZjk+CUzvvlz9wYCeDuXBwU0P0zvdWjIFVXNxqTgtBIvhPxI/LL3TLp
vO+pJNglUI1cJmAvY7pNubL/0p51Km9SGmAOtuKuGqwGKdAQRu+5Ap67GrTQquCIAnTOIa7XCnfA
zx3cUKMkw4goIu6R4BOjlWOaZqNptPbDKHm8y3etQBh31IcSvlDeZL7anyfe8qk9B6+6kjGM4nbQ
Nr9WTpQe24vCCKQXVpv0NEwvO5N3nyV46Eb74kiEF8zWdeNo+47uz68pFaVj/u26b4S+GHHvIBMC
7Ax1D4eVnaq4cJyk9oRdb6P2vkxxqoXupTKQqcdhDkHKFmi5D1LhzPwtfWwrs8h8N3yRXDcbE1T+
jcTI84xSVXVl4/xQDdeJ/xP7SKrrLJrnDFEGejAYwFu7yIn+BHSEjy8JZGivbcRj+FPsWbUc7p3N
B8dE1YFP05ahFiCBRlWXu7v3w2ZiTGgscys5HB0DtNMf6Lagr3QFS4r9gDjypu6sxglfWDE8CmyK
E5XZouHF5XE56DOzt6LWW+KfU2sSFtx9bDNDP07x6qnJzjIifB+5FUVJRh/H9y7D+lkphszsPLy8
ojVQmhkY1wnMh+YP5ZEpVwqsM+0TIkxSYLPnDDWvdznGE+nFu6Jb3rlwPSV8bQhyPVu7qd8G1A59
+aRvX+NyR5fKmoCin6EGWukghpsULV4n2aXmuSWQ6ez3j8utUDD+PjkjKrDX28h7nlyxmZ+MsBaQ
11B+kpxkHLEGrqUL0wWgtVUnj2udOB8u+x3pS+/jbOCXHIhDqO6DlCgPmdJNv8AezjI3JgfjPfbf
noAoEfbUe6Y5DrxshrBGjPfj8slb8HKbi87Qn+fTA+g0j7Q27r0A3s+PLWkzTpAngc03jEZjJGXk
Q6SRmKwjHUItEF8JKHSTqQUoV0E8kJisQFO7pWqBdsfNslIr5OiTFZsv5ZNJkVxq/vhqSUesoadN
ox1GKsZQELc5TX3T8pn7PJD5PU7OfXXMZncSAGn7kIMRTuKWXH/z+t0NPV7FPI7ZSVplla7lII+f
V1NKcWN7FEjvF1dkPkZghu9ZGvxy9VqS4StImxxQiAJ86AuBPXGRnlQOvNH93bknkDlgmBwjFvwM
SHJez2qPUNnhFLOetwOUSnOvKavMUoPZMwkcLcuJNidr9+iFoLL2O92lpP4gunL2PPZE+1XL2y55
FCOLotaHTsjJI1r9kzjrBr7meDjrmQucLgvuAqLBOKq5lNfKA2cVzvmDAjD9z+V3QrTb3Cv/RTgb
qwQqO042JrClG1IlaZUrvRBRJq6b/1Tea2tJ2VbgJXHNCO+kFI1tK+a+7Hq5ItviJmSDJ55A6AUo
mUwMoF5EvnDrsFs+Do/ekr5FcBPqmvHp6m0GzWkPIby314ieqG7VWwaQxAZuL2X7m3wjkpf1IjvJ
uX3juDSPnWBHHdT+elIrHi0LSmAz9rJ5nHL1+SbbWdMAmWetDK+QK/wRD5dSfIqS+3YTjdHNl6wk
jCdcm3yZO0QKyHBZltHA2aXKs/TSrvDNKXRfQdcuqO4aga0YkxsCsszAttwhLPvroSXLcIdxRAMY
Z79n3wa9nrqKwYi+DB/bHLhna3HEtgvm6fAGxoD33ad9Zf1pEu/yGPl55U5kCqfqsEWlsWbsKsua
a1i14L6ypzRsRkV0jNoNwWcaWdbBogdDIzhz+eKBOyH7GJUNfuraNOBRjjeIFOSc+J5GcMETRmxm
2lTQ3Cb859nBi/jvskrkgbNLjDXzsYDT1qJltyDdNoSTvlpYH+g8y74oxjPLKoasu4sObYYWuPJv
URWTfWm3ao3l4Tp9O085YyDMOhmToXBRBcKtLRV7ixalTzU872cj1ZdwZF2PevJLoFWuFrC96QRX
vM1fryq4YgmlmR8Ra0jYCqAhAWetlOVzTie1sC0S3BpHL+fwOHs9yOtXTjYx0OeTmDtBl5uexH08
d66yNxX/vSgyGb362mPXFRqoih7ryf0nLKU9TKY8u8DytMya1QNbn4/b5i5G2gv9/GBBbI5dOjX7
8+ZMQi5EF5CgvYECW4DLmKIwDYbcTb9l7RbDWeFKwtQQs4PBOgBieg+3SSK50QeNcqBj1ELGdCox
oGZMoEg4Tf94jbvw0HrY6VCbv3grBfdbnC+RhOAwxVjHBcmr53us6Rc9t1FiQ1FNDxZtl1tHKFAd
u5qmXfJHQjwPPt+7la+IH3ibZ+RdDFjpRQil8aBBty3jsxToVm5FNS8Rhz//yVvus2C5ljCZzmDl
Q1Awgf3N+7K+tLu7IFB7gKZBdotGh2nXrPZBkVsZyf8JUpP1DhdmaLD1pNN4INmI3H61Nb+Ws77y
NFKkKsRwPJHNwcXOnBVhCsDIGSD5y6rohWWCsJvcyGwP/4ViUCwwFnKw/TzzEddyl8J9tFdu/WL/
pbkdqertp5PQiR7Z/ojSf6GYKN/dTqxerzKmozMILWB1OPjv+GvHhODZEqRxxxhzHcOW9p7O/0zD
io7DbHd4VQi0PGFxldANrGbJKyEJJFa78UdzRmVNhzoRG/TCfgL9T7oki9/cTNXrvYKbjHZhI2YA
l8M+JZEJ9pZh7WOma51YZDFSGzju+IuAzu4IfPY+FmzW/AiMU4rQPcEnN5D8guZNAz3Mmd2kjWH3
9ttsBjXU+d6gPzGeJS7sX+HkalVJg9n8H93rN8r80kiIeC6WQ9XpYbNfWZZlf4lX+U5bYN7SSUME
D/0vq16C12WmWvsm9b+d3zBCf6EZJANIa9lU3zzkgP2L9WOyYifYx2be/uGzWjM6TRFql07ENxeh
Fc625x/iz2dy+8M5VgLGyG4+v1PpOsEOAaV03MuhUs6hrW95FbQaYmYuDD80VKdAxaTF+rZnrMPe
/oD1gtxH2QFv2rO5N3/te7hT/fEPbHq1dhO5h4BxLsWG5yfB5b89EdWtbXIUgBVBNIvmWg44VBJo
YYzWVZTUlGXXRJsnoIB8FUz3ChQx3spBOj+WFyUsioLjhYbBKCfz+Xa0h+1u1rNyEm1yuaeGclP/
t00ZXpa5ZUygMzckasRMkIgaWWsQbK5RG6wmtEFlSU2yiPDiv4EJg5SlKW//FlAhc0LoQhO0vkUn
rOdjpS8/gK+WE+vzE4AGB9VfRGN8YdsSmCn1nTr+W9id5tpAlI+0bnfa4rWGros0H2o66pe+eMw+
Pg3ywQzReW8CnVxzLtsM+PA74S5rIjaEot0uzAMAfCBlXznXe12nyF0V4LMg9PlmSDQXtN6rLP1D
nWXJE0TDaYe3vmoGQnd3srszEM9bxU4A0RWbhTUzbAQ4gWmvhcibL3W33x65FWd7NLGHJ3mB8m14
gXBlXd8jU7T99ssVTzHcHPF5kMZkVhlCXiu3cFb/PZV8vWxX0kbc9s0mNbFLE7Kt+klRi6H7qTHu
y+LOgje1Hj1CSJ66oCyVYUcAFWUeFHVhwVCY7WoeT9FIVneBW9LJB6UZYe3ByHJ7au0OC6IbpWJQ
yzNehfLh/8BGlJD9Lc3KiXGxWx2iA/qFYbzhvhK1CRISA1ikVi7PDg5AzwXyiQFtmNamf96sKO84
KmCy1rX1myicEQ0cSKd4kdCPWSnomtMRnVecECaPeuUdFFUUknexlDFXDFkaLLErpsQDUZA4mM41
D/0nSP8I+2pYhtW929GCySwyaOIx5v7yumaDTn1w5b+i/1hIg/4Ko/3Qf3cwTWh+GQoDJReCoGl4
xLcZbEDlDOm+GGRv54MB2WAqpzenXRNSx0PRoCwqLmsRARagrpfccCG1aOOFBDoDwK6i3v4Deqhl
JEuNevRkW2712tj3w9TDG/yv107mR5QbBMOL9HboBL5PPO/XZAjM6aiXJntVXRwkBt4GSVpW0M9H
SiJWBsEu10UEyFDzXqhhfpna7RCzuBm5rbJ40KGRx4ahZynCjDS/7Dsm0fbFi2U+5Ve5Hzt+nyV7
10afMEUPyLNoR52MG3DbOxRQq/3S8cmsGn18S1uYNBxjH8EwQ+UEcVmRwhj7D39m599l9OH4iObb
BaeoJMgcUDfitFdJ/NKcl81qKhkDewiWUhK9ecW7dEHVBvKBuxcFMf6GkTq999pfRdz/JNnNZdFv
XnHq+kAuMzzaylKsxJJHeuYG84uXg2T0XFlFK/d0v1/vFYnZu5bNrmWVEIVTfyK6ES4UElQAJZcM
9meLB2v1dvzH/y/LFPL1Ib6TibrIv00Rmx4lzV2FLl9QpvRyNfIstF1a+TmX/TT+YqmjQdy3M0B1
N2g+W2AbzOOnNEcX2lcZih0dfa+jrtRrn1hayxmB/7Ohd/JZS4avLoQGj+OJjUTWN0ODJD8UMGiR
zDUKYPcQ80ZYX+MtT8eC40cEZGXdXaTJvdbaR082FFkE1nc+0GDRVSjuFyE49BJoFFOleocRsoJj
cba4NNLk6JxrAcW6P74N2mWr5V2DOS5gWwwceWdpsfzOMtcjm1vYdrz2h8e4Rh1N6mOM4xHhVvKB
XJY6i+6bWisY3QX9Qx46xoPqB2pQjHZYYGKAqN022/5bswJB0vW45sXIrPe1rC8W2HAG56JVWwQP
K+b0mDR2FT8HW054wUmidH1d7uUN6HuvKNkCc6qXwQ6LLnuwaWzHkGNfWG0jPD1oHymRLJhPU0Ut
7GYSqAx/kX+WEnNfklkWuVTCPGCLAbViMxpF4JsHOchChGpgqexBE7ReEwCyRK7/T76hF3dPbYBI
CPZIYOh1Uhewe52mtkJim+BXvBhJn+CRhRVctWTGD73+O9+DZZRYWXEKD0Ul8VmM0/GmqUjJMSfH
ndyvsVhxiSEBPOkExaZUmTXCAH0HvHhZsX9SIa9BusH7Y1Ozjpr9OZ+/3EEzDxIYKZ1TdaB/ZxiD
37OHJF+nHdas55jjAanZpt1WTk1x96hyMd8R6wpwsKXZuVgIBDpOs6c38ZiU49kp8IQHLNl8x2dc
dI0th5gNPgtwJMjlm6UigFHtN83vahJA7kHSRuxi+2CFU0lpY72v2PxViSpB8nBVrrQsEY7mIxNZ
nr+gnRv3s/cmAl5HiSaeNv+GOc4iAic2tNuqosRRBr3xZCuZK4I1atyEHpd8U4ZtT5ogJS6jK8Dv
Z6Jx9FeYcYNafxUpYc/lx0wQjy9zYwumuPN7GSOJWrDt8mqMuangb2MS0Ves0p4wZAQbQNmM9ed1
buGsVFqpe8hdUmwn4wr1ETrL9mhcILgZwLfYI798qpWKX5ysFvG2Dwe945Os7cn+JOTY3sTSMgni
KlmfdFx/zfhRJPl+PasX01IeDZ5JpLwVWLMvdJl/3nnRZm4rh7Z6+f3W7KJLBWmKJLPt1YeVGVsS
DtBqpxdYTIYpmy8lpQ5XSC8sxliMmRBMBTGtl5PZfU0IpZkGSyYN84eUn4vuGXxBgB0nT1tLWvpD
PBfDxL3RmZkJvMAaMVjhCdEffcd1tA554Bry7ACxA0LIsP9Wh6+1hxaIWpSET0YiQF8B853Z6Pd2
O0OAd/hmwSnYBLhoGXEX8Ie+aJMpW91GkYuSi7OkC0l8BJOs2bqbSOFw3bzCS4RWCUzNxXl/B2UK
BM6P/WxbH6VnYjU4rks66CEf/TaioG+wn29nvfc80jFiE3a5R8ZWpg01+MA7tY5PkGk0amNSEc3q
wifXNqFVboZVvWdSBBJ9/1LOc/L82cSWSt7m2WMp11VMMY2zK+f/wBoIpPFIsbVaL3dFralqdPTJ
ucG59LK/wTSc9wN0esTAj8MnWlQ+BFl+blBr++XOIcsoVab0z9p2hSEnclVCXNNJjmZZabWY1JeB
QS6xBCOD0JlpuoZcIlWIqLMcQSLkYRCjsyKF4/YIeH7UKbjo2P9Wllr/32qJJENE56gSeRDcMTsE
nePZam581OuW58LwFPho5ZLc0uFy9Cle0uM8vpKHPDhJJm6lPqt1PsKdiV3ogDRNHVQu0bKHzEfl
LjuuU18H1eTw+rphMmd4saRV8C7ZhXzeOhYOU/TnsrpaMbvSgBx1GwH8hySs6k51SRGPXigHk4NL
8mDmXZl+8QSCSFWnvNZXKaI1YEq19J2fJ1BAVBK/FhhS562wINru5TSpNcSAQGgpOAxgJaS3ze1w
x8aASBhhif/DRFUZRI1RbdwePomTXD5gqBQVb10uQhcth/kbYJlUiGAgb8RDjekzS59Pz3tq4WSB
G2hQ2jIuUYdpiwCOXvf40a9tMjAo5p/+myUCCSysznAIoPk3nFk8KPjyE+2t1dr8pj9HnNTDQaks
+rjBLhCnlReVrd099jcBcNo4jUiZMfm0yDZfnOYoeabtEATZQxKrpHWq6T7g5rOeUG8MI4GXa27+
r7Fy5tUcTeGbnYe+yUEqjpP8kBmgcnGT1zqmok6M4iFNq7kO11knPbJ2l1Fx2UaAZfaNQHYONmH1
s7PlBjDsNhnS3JXAEkBsv4oPvUZ0G1FG5o+4sbIZSi1zLh5ZdRI2qi7GRQysONddxgNHLvxQDTY1
mTbGYjuSEXqiga45n2EqOISAu3gK8OBCLZJpjzYoFbiIZvmr/6zOyHP5EEJ5W7n0i8YX2Cl4Mi4m
eBDv8vgNuUyVuHl2H98FqMQc/kzTg4fg72WoxcvOgpXkQARt8NcvTK4hsUyc0/XRpgUEzSng735X
mLwSAkKKgQaVIuiT8i8xtrnMx2CwUVaXGEWDYYaXLl9wbBbTJKGLyVwG2KdLtb6dcpJ0TIqv8rq5
IX6ofnmG0gAdnpc5xr/f9vxfkiWV96+cng/JLEmfE3TKk+F3PHel4XfjV4nYc1KzMztuPERgNnjG
K7pQMB+q1X42nXZ8oOQ3EALLIgMm11/sea9MLkEWsU1T/g1btL/HH8W5gC5qDdEWW8kDvBVnC5bK
Rkm1EOrrGDi37qv87y/u8S6MW5xMSqdCbCBfFMCfa99k4LdYkJT3iIhg0WOwYwzPHXU2pIK++/6X
tiMOzfg/p7ff3DiXjOI/c0GybkkR2NwDrM5ggOUWFi0mpkiKglcZhCXwWeFoZ/7VhAgReJ+Hqa8L
tePr2Vfna+268CAHsBeA484A1QlW7bH0yUaLD7VcWMJkauKx5p/kO2H/aR7Yr7ew91C5R/AQLdnQ
wrdLRQ0rhCctqyL68ljtlRWnB/IBWTFHvS4NIJff62gyuFjMSyxGDcDtW1txoif+R7IK2Dx0FtWn
YT3SFOnmh9D8aImOb07yO64fLg5ZPN4eeHkrXFzj77oX9KnBKCQZ54WlE9GeEiwzgmURt2nL6bbh
091YFaZdOWfay+OY83lILH/xSk29Zbr7nCDoU+5a7P8HIdAFEQoDIaawPwunvBfd/tmb1T3r0MpH
lV/RILXAm0hlEg15F3i+fyq399o7hVDGwUlcYE/Oq4uGpYc3z+/mbGUqrc6l01fEcHQSF2y+OoO4
7u9aVjZxfcUZn6iC8qBM5qm5Y/7whZtz0nxFoQ3HrVcnBbdEklb8Iy/FkBTFBv1dWHKBqnLn06nO
8vTgKKH4nEFvDtj1OwegN0D0DhuyIxitnTXpJuVXBTXFa/Gg9cHsDeUCLrqos/b489RclD4sZcnU
ARYvguhWX/qIwGwd7FGXxA0CELidBbcYtkw7C9TjQbwO59obJo1ZQW19QkE+6kswTvpExV+9Fa+B
o1ftJoYIDUxDgORBqCSTOkvsrfuZQUkS9pANeiCZY7J4OVCc+zK0nNIEWiRPFiXAUNPNqJlI+7Pd
L/sLVLFxvpZbKrj1kbMdKouyJjg4sS33SIRs5yEE4Z+7VJafVb/si616MUURvOSsKXHKZOHgk5zx
h6iCaYb1d4XYQfFCK+uYY4ACSs7iSllCSNZqR3T4RmuCQkV6BaulH+9ze9fYUCgbZU/h8G9Vru8Q
n3B11KeB81TB8qA6O/DhVcXICrxsBDDaWw01h5i7DoeJt/a0e5AMXGg9vS3dN0A9s40loDJUoqus
3rI9KIUhLC67QLcC58WENi4dO/0i71qR6yS2rse4v5nWocNKmiE+rbTbO5QM1f4l6P5Pi3RG0jc0
3eWCSh65xIU4/5VBVRrB15aPrT/jIbj9bhSeCO5Q2pEYyfpsJt4QUU0JQjAqMn/Z9itG3aK5AcAz
2w6udfx5IYNaGzswRWMzcLN8/xIc+hi9okkUleICtMdpZsrbgHdwSNRhNaHvVfpRmooHsMWkIQc3
oJoyaOaSAvyWnEfoDRgDs/Cw8r8Bit9cGjHXPNnLnSbe/RiHCHXbF2WbvdjI5yS4JGIzcYAIGaVQ
0FU0senFB0K9eYsoA4aLM2hA4WnafC6L2sCQcsU4n4YG7xIqGAK5BpdutDR+c/EvZLqzgr3ptkyt
wWzyZiJv2VxcYLp5Zh7VilSaUAKPyotXFUpnIzBlZbnEy+r19mGpUV/ZbNbGh3+SXVsKOLDq6Ck9
NaA3txpyGVRmqYLj9uyA96R2+ZlIRL36I0M0+ffCNgLaLj6Gc0RJ6OmtgdmXml2T5gr7IXQlPuE/
WDA47954oBiVvg+78a1ouRAtKWdmfopnqDCGMjYHoWY/r1GyjBR1AgqS+3aaSv0wqSXIgSNs5M5X
bp9M03vIihTYw/4bT1y7HHOif5FiOlOftow8RkbVkRYK8rPlTLjpI/6Tjh7Kmbb0nWf8HvlilaA+
g7QH0ZXd8yhVybrCv52j8LofiWWDRm0quwI/fHLwUuSud13fYcqz7sgMUIAl9xgz37W/C2PEGzXa
vZfRDZFUe/GwehPgJSI/+4kBbAwXjmOnf4f9NRguA0GUy48ifOsb4VShLCJP+NPCv9nKtj+LWBmL
5+P2Gh66DIBtWKx+iojGICWiDbTLlgZa/afw6dYIcgxtsIjgxO5nkog+XgQ8GqGE9Wjee8Ibg5FO
XWUNaz/PSPEs93ubpp33GgRi86M6dOxB9BHssxQQk7EnoAD8FNfxWzxh7R415Mu5HBHKNyoTOQLK
XeN2To2LfjY+NGu2OhzoAhgt4qp8qFVdmb/Y/tZaGu587wTbqCHaknjEzAksokxV/Mm8nUNJzUzi
Gg2obMHklSvJgcoZefehb7pyxWfXomUsPibYeLrlyBfoGdVFKXW4wDG21quoulsVpFR1O2riOnQS
t9Ar25L6DBtzGjP2cj32rm/4gpIw07o4FuSYwW142CHAWoiTgWP6MrUevjht6uLTGrQrOrmEWEYw
P4GP5ngYW7akAbf151VU8Ni+6IEHA65rJ+1/zxklnybn4ohqA67jdL183EsqgQUCb5Ve9R5dJhn6
/8r1uqLP9nFV2rBpp+4Ddp9vZuVNUP1IZqYFuj9sTEPPIQKB3TX/cUHRZ2ML++H4KxxA8rx6JhNY
PgusaRTZMckZga6f2t1iqpzV0brEZw5ayqKK8+0x6P3z29Qx9FfERy3jOEqu0pJXOLMN9k43aOqb
WOB4JAVpdaUle/NZV8YR9YtYTFNLQOMcPkrtThg/dc/EvJEClzL4yIIMj9zzyRgjFdcqY7l2Knbz
Rg0wt4A8aPX5+hN3sHkAlWRNRhXc3rgUv6jp/V27NFlVeId5mVJF6VyZJ2x3Eo8qL6C/rMysJ0Bv
s2hMe/8a0rssuztEqHYjzD2tQyDoXcqDRpG6uOE39ZePj2gqN9eFHyThSWYpe67IpQ4KlwonlBT3
CNl//LqMtYN1pwrqGHOuGqWEqftMF7qOxRH1+/tp3mOAFy9iWnSo7+yFsUguB56Br9YaKgKQZgSB
WcNoHRDkMTG0bRpz1EY8sqG4nSX9zaDu6zljCrBK0oc4BGjS+xJAM9NCo9ge0EKDefIeUbbwEpKv
x2BfVk1nkfwE9mf7hLLzk7puPYc6jUNEds08qBM+2e5fIUOWz9lrq51iu2S47rnYIJDzUTmT0Hqh
kMqJxExESpfGq2x9xujuxD2kqPvfYC2AT1lRzPFerUm3fJpg1VVNA9fBK2FkGW6/sl1B8UXCrdGd
A6CYTAeIZyN30u8Rfk8NZVg0G3s2IhWH2KjtdvdOfrSePZ8aRl0rPkUKgnBr79GV7/j73wJiBDkw
sGmvDpP7DjyuEQyfemKs2Wdkns0ylzXEuCCAzyAbAKepJkMJoz0o9Ratg+RDGGU4Xi2z0kUFdN03
ij0fMbgCLbwiqd47Fy5IcaXOworEfOX9QXWBXNP0VCWLgegfyZwiDiGo310SHkUqooIQY4HMIq4c
uxZ7x3qtc2CtrDjBYHzKnQkXAKm9x8kx+0YZnw8hWMMFlPgu3Tb0PPGd6Aofg9N9I+OgeFJDtDJp
pGjTA2cD7S1zWivF1JDwOMY7yXj17rUfIhhjKK4Odo3nKBULmoAXtBdMkq2DC7dIc4JapIa1iLPr
79Jh1WOVxRSvTyuA2tz0jY/R0330n2QDlFN6eA1+glZMDt5L7KURSaUyEwZHNa09MOpThqAdYV1w
IA9zA25RwGZGlkAYcvv/Cxvm7TXHaOdeP4dma8DqgagllSkjwMsl2W62r02JY5m4bq8m0/pnwXCO
NKjmrW4+F7b5k4KP1OBW++36dpEMJlxs7sVFbJZI+t8V4dMrIFWN/Z/mm5u8GFPwM10Xs605VX8/
Qn2IQvgUbQ3g3rWAZT+Wd+N1lwmOY+IDxY8Cc/v1I3BcBZFZuC/KWwnnQdMvZKt/FBagP0Prc12l
m6Ap8nkuYhPx5+uBdQAs5vV2rXIt3NfRmLK+wXeVrHe52cNEdEfx4VDsAk1l2AsV2Ou8ukmPYcaw
jXaOyjW+kLoQST/cl58t1Mv5YrSuCspgTuMeDSfn7QDG5RhlAzNr0EwV64hxuRNSqa3PZi9wZvUu
PsyJjgaw9KItkbshD+eXcx9zglAMKlSU8RbsEaQjdFoHdK17rfgBuefXoKkohC5cF0V+A61E9Mcd
SpH36JcVsNToFzRtJb8Jlx4SY4G9EFqz7vXYnbM4bsvv2on3D44ondtAdchQRStA8uvG6p1HAoG6
k4zcm5p/4z9wBCTGTUAJwYYW7tznuyVJC0W497AQg0ReTII/dxiAcuY4gYGCltnRc8S0TSmLF70G
obDUFzFUIt+YDgeSfWP3TzVp2Xcp4w58BnrELnxMCLWp6kg9yRCIlEgQsmmr8SthnwkU49hoj4q6
zaOReDFH90nHElGuXWCi2rc/lFyHIqD/4JqYk21a++hBNqe46DwEeM1ahCvGV2oxAEOozfC/561D
WgWsYXyn0pscIvai5fFBvfsZxa826epVJ6JfoOh9iMjk1OUvmZLNXgax7xLDRpdk1hg3stscO80t
PFjO7vzeG8oxIHpFLz5ZaU3eNLj1snum0OpVALKfhFzYP4yO3gQ60GocPwKj/vOM6hRdX5L8nEeM
Zfho4qM1Agnr9wdZy6VyWHeoerrSOll9KWwp2B9LlkyUBZOjQI764WL/AWnMB7D20PkVJfir43NS
I5gSihrMr38nXr55eQQwp2OuRvef29M8PCV05RBlZnmc4qV4RjP2ZSajXLWHCu7nfrRqTCepmbdP
a4SSmFgUZkEh/5RNmI5WlH69aTFOJX03p16pssn0ofnq1FqxnSZF+mHVQaG0NWMS5+ahpzDjRX6v
m1ql5U5IaMP2D6aWzNdx8TvdArN2XB+vId/gujL4Nw1nsVZImIpHZIYKEgWk+vH5tbwlnUwF/Gz2
+h+scprwCDV4FKD+hkyAfISTirJdWUiPvWgse0IWMFaCxkDVQY4w+9Qwpqqn7lfW60TyfTKXr0IK
+JJ4CwgWVMXDRECQVcBkSrK4pFYZb61YnHcArh/lQ4Fy45yPnRrBIK0moF194D6Y3O6MPs4pTNPh
RuWsgIDErXVguVORvMpRWYXrQ34BKDXk1T7QT1Tm8ajvYq5ycTQXkIiEN8YYeotCeURXtf4cKWDT
RVA2vy9Rqf1tY82NVg/FNK1rV09adLdy65ju5Py+FhtM5zA9wUvvHdpwTZ8lxnovk4vtBo/IZ9rP
rzObLn1sZ3NOxjrJU/gBEbABowDXfl9iW3o90Ag1xCDoK/zss7o5g4skI/EoKWqsfe9qJq0y4fEI
4HaGxMIrq8ej/4IqxlRPxfPEQN2sa0ULqxXnB4Np6HDWLJxVB956H8IiSMV2hMXPbXTX8ZYtk7+U
DemNWz/uY/Q2uoL/vriiW5MrFlfk40/IA0ZzicONUuYsOMmXfjBxuGvMi8sIZxJaHfMRArqLyWZO
bE6Mf56qWwyDjXVKOXLBzrbCJ1HHzhfnfFZcPPM+M0yrTohvoalv3VVcGXoMRvyVowXzs0jd/CvO
QRQxpHPAED09fjip0GSMRqPdeL1Dj3tAi/k8NpUWWWc2ikzlx0eyQcPcsulbvVagJl3aFGltrc79
FT9sduPUS6nYCDYp/3XEceJDpOM1wDqdE4iIZZ9m6MaNppD1IqG2fNRVkP46U0GePyMu1ONfyMyz
UJzTWKRsEbtv3jVVBRPr6uZ/pRl0eCzK8XUIUXlo72qlbc+7CcwLtqlX/RQm5qdWBkFlYddtBQGr
kGAxYmijr1vrKGgwVZA796n/gaopIi/qnh6VOPj+Ihfs3hpkfoUX9xqV2lENhdS0jOGQQlrZ0erB
KmoC/na4NF9joRl2GujGXu+khXNV66cNjCDQBvMMbwsCiBNI509hY9bDe3PSUy84mqgOmCjz6xcY
6WQl5dpNrVzsB05/1NWynjAakiN6A92cyQMssFQ1d7vuyANoGOQvaf11tZ3ADRbOsIsE0LziM4Fq
nXbcSUXyA2TF4PkMPSzLkvVRgd8yzUPyo3tELQFhmIsRk+u00/bb1L352P9Y5OsQAwe2xU+tld43
SQauN5RIJ99tzg1mq3sTvW0TjQn/CZSMkJ7jNmsJ+EDG4kGbo445TSUdVWZIoENeCAY8jdhkejON
7kEE9mzDkbRX0SjnzLjs5AxiwVNAjcjV5Iz4ya3CkUdc5wfCsrUbRcGWAPwFoY/ZMSFEStXSeYOz
yQv80d4PZa338Qz/OP6StqPMUsBDcEhlwlMhLjUwAXaHwl0jljLS2orRJv9LLapiOSNtceEm+kFz
PRF+eT/BsuQDgPb3GcTR/+FMog8+9o6+ec+h8ksxoSwg94gTC1/ZjUnuW+TXN5glCWG+3mHEcGqZ
A+No6PHtJI+0yC12RGv85++IwsA08+B1Kyhytt9SxHXnS35ToT/VBEqFgGh/j0x9dTdnzzKthOlh
BS+N+bexYXOwLZs51y7RtkvSHho6ilvti0KXMkk+xUZj+rJ2MtD+gYeZAV07qovKnqy0UEnEQYYi
w2lM0UNfDenvoqR7TWMlqtZJ4nYoOy0/CgtuBWPm/rt7ALptlJxWYZ/7Dpwat4lKxCOzHSY9nWqK
bj3QVtRDeQ16JVRIuEY6WT6rvbWJ5/WCDRhUQLAglNXU5hRg7wiY1HU3mvnbprNAvc9LXyqlno77
M/jrf4CJ5aVhTJAi5lL63dBk1u421mWIAGGv4YzbkvPQHdnBnYvtWHITQzTzTiaJC7Xv5X5OWclZ
zFRThCA8qnFtSNNdCKsHTumLPhzryCglOjUVexHWeV61qWhmCEgRMoBF/FweI2sdmCFuL46hjLAg
1mOycmAr9d0zOs1CgcH00OM/JAHIsds2pYd4MPdPvGAmK5Fo8nN84FOAF3bPcQFJU4CCDcQkJFnw
2IElsXC1k4h3jTlxfv49m3lT803vL1SzThmzx/BjnFbuGtLQFTk7cjjc2BNWeL72hs68mEhysF0L
CF7Vb6MB32m8rnn8GWEDrF3C6Bh5wRTcXd1bfmLDXoNyV/4jzzNcwQXtRfNmMqE1Q0gCTnVY9bkp
14yuUUX5CBbvVkS9PTA/m7gcLoHRQSl79PgSIhMhhHEtpRW4Xt1wLh9WiOdScpzvrAS54/ZV2fT7
fjq0ECWjHGXXkoQA8SnIcmg/HZO3kbBNAqTDZUJ9dNgDq4c16hJudKLWpRJyja0mYMWAX9vADtFh
IuOKt2oBmUS6TJHxSFMgRY7qeZalqpnY+ql0kKRZ1iaJwCWkdJG5vhBz+LjrEviTnlAblzrx/26/
hRe/ju62lkb5oWKktTSzJhRg+nMbEg/o1M15c+hcOjGSetPMXdPuIOfSpjoyvf6CWtj8HqhVZBlX
ylITx/+3sv94Q8g27dP9L48ERJhAbbkl6aI9hqIWNhI1FgIAK8B/A94vQdgpsDp4bKoe0UcF4zse
RCk4Z6WPXn1p/LKy9Yk666e9o+Xbm33LayWbSTGh/f9LS93G/6hOMoUmcIh8rwgPRvPqJjwaqYmG
n+a2GcCtARVU211DLXooqL5gG2vUPUmHGOKfB2uhQnEzYxqI1GgeYCePRwLVPltnlzS/mC2h6HwF
W3piTBacWL6Ozu52NvSvkcmzyzYXqO52kmsrT/ua8FhSKo8tcSr2tHz+/Om8n4Bckmgafh9WhX4a
wevFVp6MHzsvMCwrBGPXnJYZSgeBe6sLlJt2cCjkTL3lhZIR+zlIVn0GUPERHFkiCaOZ5fzEKRuX
sd3L4UakIXN0JVL6JQy3VOmf9Ml++JJXcxUhTHNbuah+RRZrPPhuz3c9k946qOZZ2DE0PfYB8zax
WS4/XXts7K06ZHzb/6Y1SkXAhX9vAg3spOdOCj2Na4OqdxHlPMdkv1ijQLQ7gx4380kxPRuY7S90
BttzoZAc/R+JSojhEG6wD114q+rwNwJqFGTnbBxXKHkOLp3DNWTWKyK+C1OcpLFUjWtZrfaqPzpy
3NdV6GrTYc1+3aEUMxt+W+M34QBw59D7RlyEYvad2i+I/lThg/J8E3YmuqHp5/sZCRx31Tsz5LSJ
b6rXSNPJ0zX1S64fLHdQG3zG+rfSsOXNeN6GU+SCchULRhrM886xgX92RLAVwqOnhWheZqP74Sit
NVUQ9kgYt0wy8BKYakqr7+MAJTWr7u97wsD6ePScTkrzMUOZ5N8rLZvcqhm/9fdlOpcGpREFkG/r
3dvzDwiEQflukLLL+2hspQ3wZJ0CubRXsR+P8xs8Gk8Na/6CvivjnKqBZPmWZnW9n99q55RcLolI
cNwOoVC2HJAZtz3m2X3jk8lZa621wShC8f2Aza0oQySFesIDfB0lpwUH1g6/UF7u4rVpRUvPCSmE
0mVdzQzYipYHz4YpG4pIX0PkZBQMf/u6u/zNSpveX4fGwfdcWILD1olY/XpweS/felGJCFzVMTap
38rntynwFp1zCWY59P8J8rslLsg/fPYDg99eE/amNn7Pa6tJfPBmDCZMV3KARDfLSx2X93P0Ucr0
zYymQrAgL/lBh8bQB6ObaaUdFkSUJbOyKd+pDyh9YMVTKuwRIDv7z8+V4Wc90+LqeiriaGmCOEtu
+t2fDZw8zjau5T+MQkGqr4T1CYtRGJl0sp2INrVtzhnKWUaoQduvYOq4AAxbEH5MAgYDfp5VBlgy
gACpgHCDZT4uAD5c48PMiZ99+XlaYdexKy3jCxDtXgOyLK/0IM9dKvB27pkXzU67S9nGM/vNn9iN
WzQoHauoGsq8WiRsfBZqSjaSPR0YtgdlFAvj9Df/Q5ojF4VoCeo55kQ/P4TnQQXWRJhYLBLxMG9T
SSGu2eUa45Gi31VGNgV1hyHyWwniI/Z8AARiUme8309HVrJECf+galvmLfw9sUaAOF9bWN/UZQh5
6ZhBBepEPxQmdSPDWUU5RqP5SsRFbPuAFRP7j36WMOSMl8J2h86del3ba4WHnvi4VteeNmXH55xx
XYAJskvul6sSUHfYndapmhX0keZACsMEIDfqKxNNZLw97UsCaYaNr3IDCJ6bL2MC94BtAbsCUuBe
f8w+41BgRqtwp9Ox2g9zVjSGr9kfZNKWLvtdD7oHyZdYp085eEnf/Hw2XR4xk5KdyeARwCa5lzyd
iFP4itcOh3CghxtgsbluLjxIT4Uq/wiIed98gTyk77EpPZRxrCCisC2WM/p+pQx1zVegFxGUy1Xw
FuW9PK3U4POMgf/kjrPODyjiMR1y1x2ikYH9rvFet3wTrFE+rNVAUM0mLG3GOvAwck2tkGc2dDix
0Tve4CkQ7lyxzhXihsaH6C3kBBi+TT6ZsyKQ1aao2BjqXh767+Yz334E/yleT6US8t6+GfZEdlfc
tSFg7zcr56afIgwwKz15Q4gXtJ3kC9/eERhMv7FIf+oCqqCcoHT74eMdyauMtLKe06CjJYuZQSRm
5lLJ22hZ4X6YpkragKEsLqasozhiGBX+ba68gd46PhFQDGgyfc5EmY3HSKDe6IxDNLyDHZHP85/B
Ox61MA2Y5xUSTshENCtFxOX43Wr9P2tP4+ehwTcvAfu5DfU2heKZ9c9z25thSQI/DtY4QB9Bv/M9
BHKFgKdhaIozsRI/5ffhZfg44TB9/1RPiu+ewhFBPxHsrlZ52Gb/1dyC+HZavHc6p/4n+QIV4uI1
Gm0DWuNqvi3u07x2vwFgB2v0qV3rG+0s+8ZEPncEnAI/s30TX9ofKBilSx+4Um6N0eU7wncuKA/A
KNn4YfC7yimKYwzTQawsOsMh8VyZu4gjvb11wgrCGBUygb5jXCHyfrrIvWR0C4MopqGRNZmV5dtQ
zD6nVZpPnGbwALiUhB9srrytBs2fJgVjyrvZfp7nfgHTVJ989OlOb42W8ygQN/JBzOyQOw3uCycF
Sf7R+zJUpoLwZ6OXiTrgPC/GuUXQZZ76ULI8YU0ZHl3l2PY0B51NwGkT/E/+AeLhOXkKeYKIv+Z6
WE7R+nQylVi4T8iXvX+XlyOmqT3TVpa5p4Oxmxcs8eVjVaxxPe2bJg1cvFA6ZFTuAoOdOJiEi8+/
s4i92S5pfw1guW5X88NefvPiC03ry0C8FHKTm4cDkEtdiiIQVDJ+Q9k9DECMx3yPiFywJrgL1/Ya
BMsSgOnhrh+YIBS41lpMwiBoDRmiOnTmoPm6FJ2PYPE5G+aHnHH/8B2pJ3sN506dOxJfcLe/Cv15
Rj1hH52dmQ61crdQ1Rh493FMERW3xvsUvwXwAFKj7zWeo71zxylYPjwvL7kEVZwch41E3UTkl1Kg
JbPcjvm90MgilyJFSuw3zPUTu5mUFYAW6+95w3C7goSWOoabnjIEfcCenW7eewfPSr675OpMnq07
Kt7j8UjPLdmlsk32k4RJ9QWrryZ5sSBjpKI42N/B21K1bOJNv1yP8BFziVhw5UjMGZmXM4g6a/q/
UVTXzHEOSUHXbYqqg2xzUiA24KvFLGh9P7iRJ0upxc44JOQvsBQHDM8+iytDFjzOAYFxbcPZD1Cu
ZfkF4ngmaJjgdyKr4GBNPBLp/Fu2PPbPPYVs39URDbOmglF0oO0nmido0cOHcvBqLSfDmnSmZWoA
7P78add6GDxzSO8amRr/PzmPNLnoiAur+/xzxkov2NJEGcc7pmBr/aqW79iV24sBiUOb72no3qr8
kw80iXF7jrHVyZ9V8WsJIwynXEgvEiVrBZklh5jKlDrs4DgwgbcH/pgXRWUXhrmigE7/dl6JJGL7
4jpO0bF1Nif09vAmUReCjk9ZbZSGoBpJavhgnZ9sR8KVn63KpddXkSsfLKkopnO8mKzL9UKColYa
4g+J4S1FEZkmT8nAMbXWB3XLHf0xIPo4qcasn7w8SBBTokBDBnPJA3HP8gqrWSb2r9DIYn/Mq1Ua
QAwHh6xqR6qDJFUr3eoXj8P0A4+6wh2y4Pa3hpNyOOv2hpCYaqRYY65w5HpYnX1lC+eqTr6ehkQ/
snlpMJoNq/sHJPh6P+mKip9sYq8c4w3kyDBPN18zuM7EHrBiVma7O+VjZ9L87Kj3cJ3QaBdVkzZ+
yWm04h1r0mDac5H442xUagUmyeqZxWEdM3pfIowNP6T46RQ7Xh1J+0ekX+qqCUlCdh0MYhf1F62z
vShQL1MUOEp8XwCu0NlMgGR4UP4KcRju7pYQiF5Z61SInv4HmArIu+PS1yC72Y5bNE3usOdCpeVa
5ofpGMt9AscafauRi3abLfJdThj4+BF9XG/uRQj/GuY18BQcATZ2uUBlOs7HvpTllVTbQU0apzD2
QsoPqZKYD7ejgbXpYJX+6qd8qE4n8CLIDR9tNORMzYwULsVdmxkiFzNQ+VVi5B+EvL9wST1awyTx
Pps1iEXXKkfLHM9BV+48cc2MCYjwlhs5BsQML5J84kegNnebadbm/2+8dE+GFy7Rt3WQkkq3MtS8
DYt22JTHYyfmkL7UECA8bFxR7yT6py1kRxov2dFIHtzNXkyKMPedpiW88dmRqaGwtpoMBBr6iO54
QEYmzUqVqvKj8cjB9FSUTLVzJEz7qOtlOe0Xo2fNnNhxjwW2ucyc65B1FQReunKQY8TX5ZuTJXDK
hJh7YnXCqQXj5xtJ1HEtc8w1bSifUtbXh863MDGzlQZQTXQfAS5As/XqDOJWF2xKv3PdkzRCB9t5
6RXYoRvAe3Zpq7ojmth0rpAXrMLUuqOO4fWzvMB6w8F0H05vTk86ORLpFa90UTjPofrjHrrpsTuk
Vu1J4jlvTyhP0vo4DP7L+kCDbzcjCCz6gMN7gMaOyfreE9oHv25YwaCreZ9f407OMM4n5q/ZNC75
fO7cQF62DTaSTK4xrzlyXyUru5J6JCz6EvmQmFy3txrxQWh2+rk8FSA7EfpgZGJAfMwnO1mbbN+p
clZ/3FHch/RnNAWLFGXs2flsRCPhQ3MNi89B1Y59xWlgxlpyAqMYEpkRT9N+mOLBVOYfGBhSoLJw
NA1pZTjvid26WAl0s+Prws+5CpJ+uRPQqslmvO84drSmHNsJeSAfneLV+jTsI3Wym4FHT1puubQo
cfcOQ2BXHakxF5mteTAoyAEuzNgYsVyLmSlSZKLM9Jd2cWeNTY/PKoZVpibmNMkb1XU1zglAvvvD
F9LvDFO62F0Za7DlngRuyADq8yRp6At0jRY3GOc32630KHHBA4KaOi0kLAXyIjDKPtVej8kOzcFQ
7Za5J7tPq+4JOwOO1HiRTig/ggH/18etOMEsjlFd3wgqrdfcv1IELH5CTHWNswNTMRCCfhj4saro
PIbAXUsD5wG7TfZRFQfiMxVg/mksmsOr/i2LHMNEmXvPT9eYOGgSZq069b9n/pfJUVIYckn+mobP
643TL/eAuUOBDiwBmgE/+QwZXAJ4g9iNJ9WTEE07/IrPXUNqWDTDRZAjIa0kPCEQL9DpJ1LgoAs3
c2m54MQLr6PQo1Lfblfp/Um3h+CmpUqCx6aMlheVS0Tz+pR4L3FM7qHlwTagSAwYzcNrfOxz9LqR
RvJyFl9ZmlDiljZT1P0B7PsBn9l7FB+48s8xt6BbrUqay5iCUtKBmjl4UiARIOqdLK/rGfbdD+Dh
+Hhs5o/zA1U0GExtlrew89Hkktbwz9WrDUSwGZrWUTIxBngskt7Sxu3SJkhRREsYYnNi2pxDc+j2
j2Xgb1o69tDlNWWNCGzSkZn5LDcEX/qqQzOBp6AZqNJ+tEhKHUsPbZloOu8ImkgGh4CvwnrxaqnJ
r29XdLFwVdWtyExQSZyDGLdALmVQEYc9ge8Bv+MSAFpJh4SQxeBpq7vprDqUqfY9Q4NNtxliEvKn
XBaqOHbLNHjdGPlnSH5j4I4dScCH92U+1OoZE6wXlOnLziKB9zGSYj9yDq77OWMXAz7BNuvkz7Gl
mYpU4QO8ySWzbp4pSGMbWxEgt82PUAZCAFMIcJfdD1NcO5bkFQcQN6FkDIe/mrFqJsEPHperahtU
kMt2bhtY0cqxtXOIOl7A915oYNDEp5J2u3rwReiCYf4A2jEPT0ldn8hlptRpeBRyPPwU62XGCSvF
so+hFwEzpB9aVIzrQCde5ygTfAJ/rTWLSNNneA0yzo9L3/IkrrhHui1BbqVnwqHwZqLXvmpgXH63
Xw8wk2VfuYAzR8zO51l7yOP7GC3GxkCM/NpaDH/3vZGzUf7m88a84LWf6d/tkPnL6Broavf5xVTD
Kbymy1a9zLegNpXfJp8+fXeRSzqxkrcByAeqoK12Atbd4YJ2nwREPEd0hDnAgQqW43E/Tessod+a
eLiFDewQ1Mt0zmBEGJPZhiOJCGYGvXIGLSv5j4JfN7r7yE+4+xkBSEoNVGtVd4Cmy2+5v5cjp0xe
P3bobAfP91GaFILIlZibDQ7XHbjCB3vHosQeF7SmVSjh5dFypT8nbBMSXwlv6zgmO4HxVN9+MhZI
uCNCQKFktLQ10+jirbXYzBrDBezZky3hpj/B+aynptpfUaALVwYewqvh27u/XbA+2mhM6H3NdpQu
sDWE5yeTMeLWOakqI+FApAVAIAgBX/aQ5Zz2MQETMdwFpllR5bD6urLkdieRQdlAgSAYwxwkFKWC
WcEubsG97XBicohbvqvkKnDCxH/jgcmiVJpfVbTMWQYRzQTpEMzU/rIDsDnQ1vh0rzENUj5mBZtT
atVxCO3RxeAy4ojfoMI7aLWSS0BQX74EYACx1A7adb1DF2At3w7CKluHB8H0OlpdmM4skgjYVGbq
vwALlCGwLhLl9UND1wxvm6SsHHNkyhzILCUk044wxUZ7xcUffvSvXWAywbTP66nu8KheSUqYOGZx
90jGeV2USa9XdUuwf/w89XCkXdTs+5SvLEGoaoxyA9/ePiWPQXfFGvHi1UcN2dqTY+4tD6a25snY
ZPOO8YzxdfeZd3EOoZbbFGjXChIdIwmtx3FFeAv6VAwjikesI060jj7Kzdm1QsqIzfaBGNBi+gFE
PUegP/F6aUAs5L6bSmZNbdyQAJwXx25lgOIH9f6lT28bfXvj/vYGHzy32O1xO8Ci1vz0D9nAmZcK
xpHSX2nx12Vn68udoqjQaoBmB4ah9sDGTKwTo5LZYRGRlD2g5tyQ5zEqR4d4e1dNAdzrtPyOC85f
rKUBU0AoeZfzgotN9bgelQDVdNeMgvoaXv0b6+VwmslMcDOX2JSDIDswDQF76FX+3/4lrKGbUwcD
e9Zt61jnkPhYLG/74C3Z4P7hGRy7W3KVJTNR2UmIipFpn3kdbK2zfrdyar5Jko0QIaknwyii0+C2
ap9Avz9pBehTS3IFbuCCXzKuI4gBMy9t+mXK7b2CdLRjZx8hycUxbekk3iILyoPbDnxuQxS+3zuN
kXGpAoDozhYk101NQDqddbRatEpIPGWgrqRi2M2er0gPh+MWjPaVKwuH6TzlSP8e0uYh6C9EhPaq
mnQ9X+jztw89pLR+asdN1o8nmA90dsVX/isWDhf73UBLXeQ95pMnc6nYEZ/NrkBLs0LQP4UZn7M6
oG0uZX2mnaZwy/jsOyrB0R5g8mg2LtidRl1Z5okrL8sMKeRkOXRn+e/k48I6zWHfGLnCGhmgwuLp
SkB4WtDhSApx5d+9v9EzETgaufUlzbfOnXjyVYn8n9GfxRAfezAcYmOscZSIuPcztibbwS4tO+qm
3D7imJKLbpxaT1nSC9pmAGbqYtPvk1gwgwdg9D9AQZ2tRAsFhisSnHVX8JOg2JpcHAAzxMDM2nfQ
md8klUNdFk9o7Y8Sax+nidxy0/+coykpaX43Se/7efwCOhLti+mpGjs2xcCNh/fpqX9NoBRyAXma
x6oCc04/uuFpFha9l0zjB7oTGKXwhq0ww9MNAjK3rOYPEv11Nyuq1v//7grTb6oP87R/sJWlByLV
JciHcowmR5IvlUQd3r99h6uLYyikxq5P3tgf48YcQ9Kq8i75lCU6RiTtp9yNVbDVah4wI9SL4Nn+
cUuEOISzsOMEbRm3GtCa0l+XpT1sRmD0Wsv12Z1g08MYZAZBjzWxbDk32iIyQBGpD40sc3ozyQ58
g2Nhc5ON+xBJ2pOL8zp+claMVIlH1AoX8jlqMCGZGu4/FvPQpYfGGn8AbKugBg9yHz203+e95e1u
VdzpVNI+ZMeYHiwoLeJWRGuKjMyIfgACxtEGZHC3nIWFik7IZ3yYAU9QEk1t6aN7hJwY8u35STpx
wIU7vsSq7WYUYcF5SrhVpajYUUcSMcVkVQlehF3K9K2ZKOBjiagKm3Z6n+Qv0cmyADzoh9okb+iI
ah4P9MPZa9iZwlw7M6pNHlVy/7bJxoR1m4VSumtW31C4AkLUEMhrd50IOWi9jCUivffhjAwxmPsH
21GbiriBepX2LikLCasp3Jv7OHxzGKP842oSVq7USsdXtQO0eqypi0sV1LqSYq830iIdCUFgTMDN
t6xahxJinSEnFxJVNaMUCgl92jbNtOQ/U16ui6X/hF7lBH9o0GbgtFFppWiTPs1keI0U4AEzYLmb
2R0pwFtBv3DWhMzcgNcmUkWpA5il+vESqWyYCulAhIEhYM+LbPIfu6nS+TiRe69IsIQrnzTSBdz+
+/S8K/cVqXm8lx7blFD72XGlxc5+6AsDNYl5iR039cm52nfXAwHpoNfiQCAssyrpP+IZWwEbl8JQ
b4L5rvF8SvPVs42rnsG6EmFVbrJVmz7+agWQsZo64V7ZaXuO1Ko+PQPclJfwOwlPeU5mbI4JSvMP
rLcPecq2rds4TznotJD12AyIajuMws4VIOYxYT7HIJ+SdzCXFNqRzSsr9oQkHqXEx7z63lHPj5GD
fSnLZS3aRnqj4aEV2DXdTZkfz074/BA0aZpW3cUw2uhysKN75fE5m0fsC0jMHqjtw/WVtcSzz+Ec
XS54vLr4c+bfBJh/khmQiojY9yt99rxA6flqKpkS4aOtAOhF5JWpKq+AvhsZ251nHCgRgXgPeqWg
/xMsxjUVQAuf3trby4IDcYpc0N809xUMQHynsDtAvjfEOxUYkH9S1oXS1yOC73nSG8710aT/TxSt
01fKTNlNHa7buG+ZcJ3c0OmWs4yjyb2loHzdWXbX1Ll6BQHozPs2sQkWLSepoP63a7BhfHApjPWU
f92hSkTTeR0l33S5iwrGGqtvvJ+d9Qceow0eVW4rPz87qmyl5p7omMTdFegwI4E/yp5ykk01YOp8
KN54tHNPl3PmgkdJMRVIDUcYdX4shp4kdUmK8vqa6zMzdoEYXl97WdBaP6G41+jrI9J4ni6EQ5sI
6YdW1D388R7OlcCd9/Y/v1FyBhNISL7AbOlvcZwdpGOkQqTrluD3LGtZX3tnaBdbN0onIP7xZktN
VjXboZ2x7NT898OT7eNQE/txziPUt5SvPl6sAYrknfuqfIJmL4c8pfbMVVWJOzrza+ln9m+Yh/bn
uigJPwN/xbE4xFhIHqJ8E3UX7gW6RAl97WR8KOVsped4z7PJRQfLGWZXJJkqw+/MdPjIne/V9Q4K
UlUG8EyKldifUi4pKfUULrjizacmy9q2AcgYD68sQSpoRBiU+ENsaco65J8eKrXUaWWcpB1s3SHx
RygzBCJB7YgDRCQAnDDOkYn4CBKnYSXzu8ubrcLjxXOjv0rcaxnW2w4uCpXH2Af4LTyENt3ZIv4f
jasE5Fq3diz0iXTPlVs1HSv41rUE7XTBigp5dx9PECHsUu4iKL6LKXMGuXHk46x/9hno5N914Jgb
3piT6ME/S/K0MngcFybhoPBYbYYABKOEvNcalswQu7ngCrsGboWsMbF5Zn+5He32j+gwJd5T2CLJ
YL7OKT2cZ3FV5wK+Z5Pfi4D6K0Ev1gg6rmn5Z0+Mv5WF3qRKHddFa4OWVz655PF0YphBU1gwoPhc
LvDWvdSzn7pqSi0+owQtvKSrP+a5ZX0aUQP557sY6MYf1t1LVfVN5dcAXKHPUMmw4OLplX8eQEuI
XU65qr0+4io06DwJsiVoTVSfII1TW5hyBv1wJ/SE32PyUftvswzjApEpAGkq7/kBA0PMYVNqLd4h
OtBqGRv7Fl0GQITXWaWw+KjaBq9F9SSCPGMRylsaxl0epGJMGlqRhFU5bc8DD6X9Y8IlAbpaNJK1
GP72sK9Fhzr64QtKJ0ZTyZ8gdTqVp8rn1Iwe/h00WM1Mt2+6+RlHmocQ4HmWMeQWNToz+STgZaW9
TBKjWaKRSs6x+lZc7XQ3uG+D5393Y/RWry9xLcpVYo9ctzMFEEEMFzXCD70SJ64qCHn7tM1c28ES
m6/QDX7Xf6imHbUuF53fSEWGn6qiCrcA6sbOBc1S01zMdh0hzjB1MZYS8tIj0Y6mNK9TV7H/HvZr
Yz2R4qq4RN9V6Cqq1UNsZ3pUx4BlWOzTYnoUp6HclMomm1nLenzy/TddEl+E5O5L9s5b4TFqFi1a
ZLdvEUy8tWIMtMwgTyWM+ZaKFQQhYnhMfreNHh3c968WLLBWMm6bnFMmoqzbl07CbMRv7bovIZdI
ikox+HnWvOA4pBgnhwMrNRPcOLqkTMEvTFmUmheCDtNaMOSaZ3CRwrT55pxvkpEBBY0+d+9I4VLa
6zOTLELbz1Ig4AW+P7evcW4DdUIDSJWQFXE5X/tCDovevqzjxAWFrXw4lgJHv2GpJFO+Wximr7oE
QWewqOuJvcag29bS4AY9LOZjQztJrnvzKLlNzf+zEzS4nMK/6v1wbub2MThoDc/VbFx+zlZttjNj
DPjhS4Coo4xsxYNuWkBJy4IHy0PHsU/lWlGYtPcMoef8Ua0famuXI9cqtDWp25tuFjwJmaTohiNM
C93JptvAk1Smefw6+EY/r8v6WV7zKqXxt24ThjQReMtqMsUL9VF+V5SjCmO1zcCMEOe9YYMLb4dz
CveS31bwqMEbin2zJVE2jC3HmvjEXfCjog+X9BlAHMjJcE9f+B5NQUgLUIGFgKclGq2Po/zBpyz0
KVRN8E5RWa38oYfKOtwH6mfjtBxn8rMDtDlLmJrhmxqh0PT6mFPod8+a2jp2k4bMgPNBXY5b+2S0
zGs9YLzKvjAL4eJ9AR+0aAe1Qq/Dnk4iowEIzak3EVSFkeZ3IpvmxOF/+2bv6HsnzXdsRPA7i2jR
qIagZ3QMEl+Zj1107jFnl7UTkqbUxE3htxU8TFZ18pujyX3HsdmjPErO/rDu4GZhi68el1cm+2Jo
cnkkVqeMSWUyWWmlYeVXkuAO8sWtAawVFH6i9wJ1HvAIz9kkNCsnRhG+6Y06FvUMRW+UqN1WZlQm
RerA8+LL163mIfCgGe7uWbZvhihonzLY0sGg35xq0v4yYcV3uv+g3Rvk+HYBvMB5/OKqm8EIZ5Ih
2LyZ04CAKsMdgghVvmtAgspSBiyiozO1QA5TjbCMISVkk2l1weUmlmnnFd9JJiRQ1NmE5jVXSvpx
AvSlBfoHcpaPs3ifvVDMjTv4YGyI4LILfli8BtRUp/KUcilojyyT7qMBROvimZnB7sSdohKwmILR
iFsWTUIRKeyuduwAOwRqehIKDAGmpRudR/ePc3/tR6bEA+7XM6+qjypj9doD8zvSabtp2cqjwpmQ
IYWDrVQov5lcFEv+fDlIlXc8sIEdVRz2WcKl3bgYWL3vLvqKn7Ha9a4OxoTF/fy+SnVkin4XoQfX
ss2Kz8K95Egkp2pweBariGYTLEvCwQRYplMnPTZIc95kVJ/RXmNECH8u+ygZP37fX2ihPQvVC3oH
Cl9IhhB2wE66l/8IPyjYox6H2D1yvIoJWW7qMdFq2a4d8W+NyYDaTrHxTuhblHTXeBEafJCrPNlt
y18xXCgYcef7rQgQA+S5tGFf7PDNjDvts+mRjM+9DLD9k/kMMa6/IhYSkcom9GMWhOVaFYuTHRJq
QsnxZE7WUOFe6L7Jeb5MQ3wstIaakoh23s3FK53U6NaF5Y78aa05wkJciNhFO8BT32t4OWY25t5t
MEdg/g2TTkv0emNfnLG13MeKgSNFuIZNdy0pTca+ca1WpVYVsW6LFn4vWzR9zbgXiStO7zKYitxd
4Uf0rCZ/9RRUEp0RKI9hmBX0DtFB2u7nBovZBoQWY+iCZBgDhf2apoIPQFKzg6Uoc+krJct3wYo2
O91+WvI5ARDEpFiiXq62KwqKFQfRBwaPT0dMadpJQ0IUE2pGNvRVdyIWMKtf46ckSjDqhF2MbkaM
U/nXsAqzFWEtT7l3U6O14l92dKL5E5f/PJ4JY/6GCC8nDpu3o8n+Xk3JwXtDOdjHvoyyhKHnQexh
v3I+rWLyv08Wyqwqu9aelB/xwmRFHtVcmWQofytg2hqo+cXeS3bRTScz58xFgPc0T5RGDPxH6D6/
c1Lf2r+lE1noRWxAhknine2mCOQ0D6hCQhQopuGxl79FHI6HfjwcKulA13uzYRfcHA2geaq1j5WU
b1fCFJ7esocZ+Amca0eXPBjc2dTLKaCySk4QQO1mET6PXwNda3ZkO4BE6cPjhWlzwSqKHKPKhlo5
Q+60ly1Gixh0kj0ZK27uFp2Crhrns3LWlZK7eUiog0OApRYMI83EK4k3Feow5muGuLOq8kwg9XeC
qVEXO9L4fn/nV8+j9hVSXacAyVAp9V0JX6DFtDuEDj5oSkulWL+I+xh1Nlh6kBTjbR4YL+iqDVx5
9Y2Ft1yqeS4OSlnLqWQDtqULQmaOy/imdRacLtwKOkxKJZoFXvoaMAgnQzJ2VGX1bj1YB96ygJ2e
WZBk7pmNQmbQ5IlFzyl0Z7gDIXqby4csE+Jj/6Nf2l6dvbqh+xCnuWFM/GvL91KFc1roJ4NK7MGj
hx844TADp0guFIicI3PKr/XyuItjJ/slymaSP2BTXiFE64jpUO9SdlkNr439WgDp9/tmL3a3TZfL
t5FlEPzZzAaZC5QmYbOaLStLhL1RBRJMktgcfBpE1Dlq4g/1uj/7nQQVYS0PIbzKfPeiqTot+MkY
835kLWl5Mes6OxYcztdRhpb1/SPyuO3kc1ei0qGCkCOYDOE+9UuT7G9QX9uBlAe5TxXdqHhdmeyp
RGLxOJBGH4IO2KSLjfMrN10eh49RQ4OxS5kXuCtl7W8vhHJk9o5ENd/0MyjAxbYZpaI1GsssOi+8
Da15Fyus0P9m0lf4VfnY3fkLsQj2CK/jrTjuwKdsKpmBaygfzo7k/vYNJOpd8yzFOIWNgR+ZGA2E
CbkEj3DUTy3NLd09R/P8VKnEmgVgibhpDGZ5DDCBkdmo8KqVBF790FiJL/yz2nOHZbnyuDjwkd1u
GY0/EsF2tr8vhJCE+LaVhxMDZfxDPDZYKNGjitO9elLwCr/BbiueWY/qCukqb0FjlAPcpFKozo2g
cyqZTM8VlfVRlf8JfhXkbaXMiVMvkYR8fz+w7IHnO+uxSWFJDa8/+9WEWMRUTWGbbpaCxfF0sU0i
kimgqLvHdpXbhJxz46HEnCjMK2MYYpwVfaBJpUXZAEhRf0bUWL3viLctU/lFODsrUR9xD5WH+Ioq
xdqztdkAt2GU01k3m+c7n5waq0V6MmNzTrHnMFJEhttbYn2i92ejVCcDn632cpso1AcYx/fe6jdd
775oMwr1U37UErZg0iXHLrMyvSQqRXbwbWiGx+Hv2tP73aNSTaIM5UUwMsfNOm6OWb9Z2tqFHwpr
0i2HZOGo6l1f6yeVBoTl9NdqClLYuNkdIBcRXl6bK6VuyaD7YYjQF3ew3P/5LSJYrTByvfp8IpgN
WZCZcC1HqLTouXXF6BLcZv2aO8cuJoRqC5TaL6qYmv9hkoT17jB7S3oUFIDjAMWarP19U8e3CTtW
THtg9dPX2wCTj16p1HnCQtCRun0gJhMeVbNAV25ZfGy7Ih8lc51SwC8rFJLiV1MqP21y0bynYy6F
m2x+S47unG7DoqigwZA++Hz7xdStSGgDK5JjNRq4ON0C2OehASRXg6DL+Fxc3qXto5/AfPhV4cud
DeHzBT8pSjt3DfN9gll7qNZCkGMCQ70jRzriQ+9xSIqFmeKhq/MeVJL19sMBXPwc+BWx+6eWHppu
Hx3texYeqGffP45GIxHzAl/pJwm8YwUPZpMUJzpJ305K/0/CQJsuNQTjqiuFFO+eX5rWr8U45czY
nzBFYVrNKHAULZWUfNxg3jcPgA/vhYtZEo372CgnY+B3IQjY6nw3pPuL8+7czEnPiWZT24bu5k28
5zB3346udQL7CTcLet4GUhRl+ugT8DymlKro8pyKaCqg1OBtk86nkEYbhYOepoTL3GdpZNenYf3j
/3MNOlc8Gn1gr8gjlF7FB0kcSqBVWCF0o4UMdq2rUqmMV8XDdDg+wFCEWZy8YllRJSgDJZL1KK1q
x5Pkg1gkGXFzui9BpKIou+PGIyva2TANqvQG5sD/EQhzsGs1i5FQrE0aGNsZlnODVNgjg9FU63r4
i8lovePzhCo0kicqqy5mRgMVY3AEODQGoePjUa2wwAsS85NhsY41ytdM/qYoVFLDqOGGztM3OCGQ
0bGkEMnZOSjcgqQIyZC7ehXS7SUmwRVjIErn/zCsM3NAIsG8NYy6nUe3iKS6bVvvqPz8dR2ST9qX
QBnmK53S6Plc2WzRs8O5HLk74leyYjDY/1OtDYTzHsmowlCcOQrzZj0A4f/TliofBuV5ckfiDATx
JQtZotU+2NNTx8LgyV+4GY/C8ncMYCvjnlf6szfTWfyL44f0zLT5nzWXIYjiRB2mAY1UmniER4jj
pZ9h7luwVdXgHzUUo1iCl5v8sJtYsGW8Z0c14h67qoOb6hgGzQ7KaUpQok8jsNfZ+YT982CIBLnp
ZDJA+nmWPg2kzOPsmTcAEX8Z58wf979PQMTC4oGqpSH1n32XDYGDKp9gM+rWRhHG753QJuvuaYl6
GZeZwg5gC0g0fbFsgi2giRhjXpVhT1EcJNtAoP/s9AHkXls/R3+MguChvvJzQp8D5vmnfoK237/s
bp1wp3gRk28n0cmovjjxdndy1lysRW1qZKrb69iVoDHh9JNE7gdxRfk2ZqnEuJSilUfZXShgO4Ad
RP4LuXam0hfV4nII+TRwy5UFeMEfYSH0ByvlVR7Bpz0dizW8spgyBeguXSFUgN5AMSjrs22utCWW
dTH9UUcskktVyM8NzkvFD/6bxTH0poDb38jB99DHTBGEcbImcHcWU4pBk5Hs6sb0WQTxYvY+mMR3
PJBkfi5It2uSpnKSrFc0HmfONXODu15UHhdNyos/OanfgzEuLHPuWzdH3nS6Aj9T9A1OdESOf5AY
6BTunK8ba349CjcLhKoj9DK3kZVDayJYjBzWb8n4ZyOAwoafVxfKUzVw25cUULgtdOJXEVDmkk85
iXCByPMMVmDN0v/5mL66079DIc9KB9yQYfdaHMgElMVgSIpTCEYuwv+iagHS8E9hMshUeFlR3bUy
aNi3njUw2cp9K5VlGO1aJjKVWMrbUDdwag/UDK+VguS4EvuMyIuxvXFKQwxaVirHKhP5VOxaBFGq
YMHLIbeXeCcsrRSWG8UNu6uNlh2Wh/p5hGOdQ1x7UjCoslbGJFYpL1zr+6XOJHYDEreXdnQfsVb3
6iSE2THNYoAx5fgfCHl7fOFcRJ+Y/IeJZhpewOTjPQRjTZ29Yz6DyMaEcARZvFFqChMkyxpRp9NY
ogPKXMsisDok5+XZcE7QhgizfKk2egUJXGhlZlR7ThrteE0GNTvGwMhzJm6HdX78Wd5z9zxpzriI
fmV/ukwtsP/WCora1DUZIj+n2tw1XzbMLLubPw9LSdldq/YmRqnj+Lklv+O09Ska3uw8MzI6LGWG
4+keheDEuGqNfuOiHRhq2FYMcCbg29rK5N43aH6gz7kGeOYMfeGiJ7OugE+gl8Kn/sEIUmEE5/uw
0vLYego7m9a8sVISIH2DBAW+v4swfES8qgwz8uidD/MoptQ5BR3x2u/zF7Moldr0107wslAAW4Wj
9O+SqU+NNKhWM1fuqQFO9ZBQHSKvNIaV4tIcis+QXmu5JVhtUTOvsRtHcYs2fXiKjXwDTtc1iuyw
KRQpq36w+DY572EP/J7q1I6gu6EI0uuYG+rqxfWfXTGB9gERXSGn8sAKnbZRP2JvykfsBEkbgjqt
+/9QVa1qgiyerS+OXz78oQkcGiKKw7X8IRhtvLZO1eo2xCQtp0yRv71UhGky2MuT0x6uzUQagmKf
7HUKBuVByoX+UDNaeUw8iC8BMCzBiVwy/WpDf/hE057YZ57woY0ccT4Rg90Rm2G+8Tm0mjQqrcZc
wEXF0qLbOQcW8uIu4jNcfKsfOmZZGfpAsDDYVlrOBvdCDuAldsXLHTCVsIbZbRQyJ6Pksa6YcheM
Fow+46EqmUxqtckViv3WoKw49gDjgtxWlLs5/Lq5FVHadcJbmgIVunOD5NaOJV8sGawHThxCe0T3
gZGki+FUqJN9OMOk0u9jOY5JLGAQ2priAOso2sEIjfD7lWGZMsw/3ExryxbVEopC3+CjmSYun2Xp
sj7r/m5QYMfNOf3tYR7pdnKpw2O0m1LZVmxMtPJsNlT1AI8nBcsQ980x/26+BHIKOtX3zlcXteUO
D4+WaHwEo1w50z3oH+lJGAoQPc2KRA5sKnrjw+SkPilHDJ2eSup18pCdqd+/BO4ck+srusvKrwBI
DPMVRDPqd3KK1ZXnoA8Aw6F1xOhDG4Wxbf4wbB+1DceE+QV1Kn0nb7EcIpAXPGy1lsFHjihuSXl9
m0g8I87+9fgAot0moGzRZuLu3DJW4r2eB5Mews8gl5ljoPb8unoVfX9u2S9k7+tsbpVg3jDILsF6
C+tyNKUCAl05m3GE6wNNsL06C8hhuQ4pxL4dP+UzOQb6+ujXKAjm6xhpHZ2Ul+I2gAvoDXdXSmcA
9iS8gQ8R7S+jMXfjbY21C1BIJlS+c2xZ5zpa/LTMiCn1q3Z8MzH/Z+hEpr9YDe/WAnyl3u5o3cjX
p5KRWcaXgZgt0b8muWZoKtxa+3KRERPzwrND21gjACG4Jcf9bs89WAQ2Jz5eICgJKsRVBVcZOyvr
HzoyE7aQ6eDB5r2+2JN1AknwYR9HgxNekRvRgU3u0ZndXEYfKBynegU35FSIOwTd8wkCxPVSScgC
+/YC3EfAZxmIVXjYAjorLOWPafuCNlL14YlkyjObFRmMfbQdgJVjrU5dpoJFc9y7gdtDt6+E2apC
BL/PzLQpcEfgBjhOzNIlLyXbtcfultDACX41TAb/9VpjSngA610dzo9Q4teY1UKzLOdj4SukBzIL
r03eWYMQuOKW4WscAxHJ/eMLBGkXi+DE441spZMseqjujYKnny8mHsJKCzvNOBneipLU/safe3XQ
JoGDhx7hEqhh6Te/vs5oOXz901BR0mbcBUzXlo4YJqPNKzucX2n6cif0NAhn59RHdW2zOxWBLk7W
RuTtsWnq1vaxTuteqkr3qV9kGGMXJs1gO4Pxjwcn74TRFVObQ9zb+JlL8s40LtCC1a+MnTOYMUdX
K0mCv8UInu8xx+dWDCayhUc3/BPhxHr0W9t8Rra95MTZbspyMSKv9doWer7HOUe2OCvt4rzm5wHf
9QQCjDeIOGCfogleftB5Wc6WmiBtyYHQsn8z1EEKr4c2OrYoq3d02liVeQVd4pryBmAWIePx3dob
RShdK9Q3tgvxWdzQ8aZhuYfNcHziA5WT+y1mLvKrfzXiI4YnGNEF1ROT+3UpxwAOc+JFVHIt2Eko
gObloU0+2BW3jGYsL3h72xvW2S1ETmftAqOdxudGTvd0ROxXHSVVe6TW0DQT1Hq7MvDVsr/7qtCB
DE3+QtBUGfQrgfImeY3Pkmf/p9962uiCRmEreh9JzqxFeoECRr/jdB7NPIU6zTg8ZgsZl2tofyQV
7Ai7vOQZjtLOix5+OuR0USIcfszW0rbmqEQR2CtXH+AQOaYoMSnLg/i+ae8kha+zdwrWLbNK5LkF
q4o8xSafY2BQrVfkH5qvGOLFL0VT9o4NePor2pY70tH035zxf3jFzumqzPpkItZZxa1bPpwykhz6
0cLzFMq37qeznHfOhQ0n6LFTP5QgphfWXlsVe8WDslEgplxSWu+LPuotty8G7x877vaScTngK+VR
BwoAQK72VPL+8iHJ7RRH1XjubDI5vp9leP3DggybaYBYRKMHfSEusa212KWoMjJ3q4FFPCdiEhAl
7I2Xai4rhBANcSBn0d7RkhGGSOT1EiqRwxbwPRTG1zcKQqnlZJOUuac0c9UmtoX2xu11XRrrUV/J
0UWZ0CWGn87jTTz/A43hdw7+RJ2Hxp8Q9C+Z+uSDOEoXVwkU37DEXz+BrwUPTdc2CEht5+D5FbZS
NpqmMIBMsRorsBIId4rM9ZdbDVU/SNSCbwJ9AY5VoTUH8NPJ6Ns4iGluux6DTvy9YsZDcWw7Lbsc
Xj7tH91zwukgggdz4pP5+8PAFROcm81Uk2BVgSoMMOXKyX8kOJD9PFawZY+pJMIjUGGpCv/fkzy+
SbvDR24Znsz97gI9sXHHf7ELqV/wZYnE8H0ZepqzHMeytlw3m8YHkX8d34Q23H4VGppVjgY28gjT
fdtXNzMWp86uZH4ZX7W1EgYJBJ67aweHHX0DFdLMCAvg/ENoP/0B6FjS2QSu/B9atoVT6B9JFTZl
MrNDdHGNlHoz2zp4AjvPXRRBYj/a/a0gZoS7E4wdjY9mHBlW3e/0cO31HhKJ7V4hDP8+YI40Z1i/
qOuaBTlfqMTyMwaVSFQbXLD6X2bQws1CS0+0aE4JqXMav45K+Ja5l+f4metaXLG841km+tiS49Ac
2AMApv196e2KTCTWeUeXyh3xJn2LlVs6jlPymKpV3gChf98iuegT4+6tVi+LZ7BL+c7eHHXTjhsQ
eDf3HxsRPZhRvWQ1VHqJAjULE7TELc5aK6R5A0N/5kSWgUJkJe+cvXWjgy+8IhdlIXHN47UrdsvV
FfhzQTqSwdkm//mr3la3BaOeG5tL+QfOxfHsqvd6ixiv4G++QCpXALVBaIv2dcG8Y6LSORN8UmMF
ike4epeJn6xWfHZgl4rHh7hk09WOcyq3qb2FWPeMAkOo+TYVW5RHTSi3gGnpq9zoCBkDv22qmGLW
mOZq2XbG2eLN/o/iM4nijjyogaRkhhlYwjMSII6Bx5iwQ2spsc/CU8OvlkgYn5IHgsEkh0G0M4nc
4tiWouTE01X4NeEaAIFwMohyBRK2U6jP61uiQPGyx+A+/TW9i3BsZrvdGaQjwdW7ydTQ+OU0jmn/
403BRMxLsU7C5NqI1lpaELQdeNVqe97ItiJSkVOq75XgNx1OPl+hyySOPDBIJNed+XQlwpASw+9f
gJzhAq68O+zJz/DmOpT6B/4kKGRE3hYUJGjaBMERyLzGSgEdsuYrtpgwZzPQgHV8++Vq/scyXNT8
M+tEMzaJ/+LMpgxzwQEgtL68QNYCvK3E5SzGPugPChOrzyew98FWJYFuSXJdGNhZ/a00fN1uVkf8
TS1IkfTOYaII2UVaeGM0LQukj9KNvp1Sy5vbcG2Ial7iRTrFYP3VZXFpoWKhMtC+dNVV9UXYqKL9
Gw3zu3s8hMPFOdawWA/xHr3Jwgao/7RXhdejYMygzlFQOKcYbtV71j4RQVx6vNmauVSXyWdV1Q4f
mJ5r4Ou8NFtsboivdYIKhL+1RLcYTV1LILPuXVV3We6v+2IuTQv3Wi9Y09QYquGoWmb4xMFH0cjt
PsQUCvaNVWGuA3N5CXtHFnd98CQzjxflmjmq19HSTojvtUeRDSkAPzlrNdItXbaUqSTRBVCAk8qe
/6EKJAVIfmId2oub++lfgHFrzieI+dcQlozLwG7WQDJiulAKHMU9xp/hUEECX74sQcO9GzRH5LaP
uJB5y05QGw/SU0fuRWRdZjx/zZ/dH5KAXBPq9J/YqbL/q5PnEZP5fWdrGi3pyKvuY+g6sgPKaD4A
/QJobsX7hPBj989z5KM/khbr1AnVTJCgFIXQWHv6MZF7ZInxdDppncDsic+EUtDvxDqMaayemtT5
m789SfuT8hBY567jbBFVSTK37MFV/lh9Og9U3+LitCChQ9PKOZecyhdOs7q7fIAklQ3ypwocpPGj
IMTLCMZSANU/ODnUMJI5GAnpPzkjWTJaZBrIyU1iwMB/OzBxlVZoS8sD7XbOaAh1TeRX8SYN2x/u
YbyakQUAikuimxVICgXxSeUn/4bYjI/Zf+nTdy0j9UWIeb3BfYQab3kamjqmKBYWEHbUoUP9JckH
PiWv+1P7dsuroMEK3IJ7PZiOUpPO2hTR0AbBSccRqW2zl/Ite4YifyJIlJzgcnlHd4FLUQY00lCH
jz05qlQrPD3etOOldAG4SGqcVIdv+Gu/iHEw1GnhJj5Qg+sIU9HDY8BSmJRzN6edzy85BoUD05Ob
Im+3IT+leaj8obXn6sdldlrXjyCFYI+gE+K17JkhoS31F+DwN7dl/vA8dXf76V5TBxnmWS/RiXLQ
xqxiMmjL4IhEiEZGSyLdoQAMMCyJtSWvUDLJ/7o/03iKM2EZw0GkAYqu9N7R43D5vj8kCjEB71PO
Y4Uqsa2QkF86AabcbLERvucLKMQRgD7WVQTxermAmNxOQJyTglqcxYuwmeAC5sR6IYEcdPrZr8BF
Y+yuFu4X8uBi8YxrM+6VM4XSZ6nBISPn4oOomxIo5QR2/o6oWV5TDQqW2iSXJZf76rKV2MwjCZ5L
VW1qWqpuAzM3FKIfejFWi7rXJykDSX0puBUU1UOqrxPT0WcSBEcAivjdBcizGRyAXwAUB7qgHJm3
CT2d4HJhNbn0O6esDPh8pLXUdsp5lYxlxNqmbsL3KQBdExkKDBDsvlBZLwMG71CvRfH5EmKIOMVs
65tSm4aqodG65mefTN/T7gBcy0f6D/YYSfyQY3/8xNBfZR4uby5QA/dlkIPBypjoX1uVCADdyjbh
tganprV/GeSsZ/vT9wU/VyIGzP0AAcS5/jkvvvR+aIEjHP+JbL+Dpy6PSnygP/Ple3tZVvYVRacl
IwZbcc/vv1QBBEj/B5j+Vzl0okxKcHK/5PXOiqlu16ZroN1tZnZAQ36VY+ZwXZnUtGcTFWIC9kq/
PdPGmzPpC7ArhkjDCGtPxOIwoq8GrPuqO2Yeb6/L5Lyc+qp5S+l/S4J0wtxSW8HZ7a1+WrTHYxX4
IDg43ZmNv+Zn7ZaiqsUnUBdqly1GqzCxGEfX7hSKhVdO4icx77I+xuvzcYyLFlFSt1j2pcuxWat9
U15vOHY+DJfcXqHfgUSQy3UG3cQojAvCdIew/kHpAF4BAb3ETngJoKukv1mkJZN2mD7Z6I4Lh2iN
q3EjswnYofMJh4mHUSA4pEyHecp4DZRb3x6IFaHNgJ3lBY00tQW+9ju72VNqfqnJtx3WH8uSYxkI
uIFa8OGTkmH5SAZkIc4FAWcox49ZhBt5sPBKcwizVLKRAgRTIaMLhgvzFKRjaYCPzh+WW8YxvVpU
lYg/5W9Lga0s5OuxQrImuF70i+4ihAPtIiJ2Rd1c7ysAdNl8jwkCY5Q+GL2sgSfnUU06Xi6IRr5G
umfF7lfTw4eMZ97EJTY6a45/YW09IwBoNlX7YiSt2Y2wHycos73NIrr96QmYq+hvi7JKdQEMODnS
FPDrTj+MK5S4kuPGG3Er6X3hYqV5VyVw9MzVqk9u6i20wH6Mzeebie/KCk1OaUDf6VLc6miTVVoo
019yCduqtb3sD2lZ1ctEEsJYnqDU5WAyF1XwdHTURYkpMm07QGm9nPm0P9/T4mymxDAZIAmMYS0F
5txJ7qzWQ6KLEJmuiXNToCUoJbp8JVbBEoZMTSEfDWlgxr7CKZMhgh4HJbuSZS/e8zZl3uT4R5jU
PRp5lrNAP8yUG3+2uS1WhPvDNZrtM7sioD3TF2UbEQkrqsJXkYMgXaho9PvzJ4Wt4INbEzagFyDY
txw0WWgnUFKPKtS7LrbazZBsK/z+nBiZlHUXO+6EkP5iPAgFUwSfioFrScMRMkCi9SGDCxCgicil
mM7CmKQEwQJrD2OCwy/2ZTZS2HUWBfouHCtro2ss3X4rf8NY5mciUbWKqVGBONz1pcQThEh3PSHV
0Ce8CDKQdQbi7YCirlO03mknkfJxFA0ep4sKc9DaOCLdQvePFVyNxo6ZSK56JQ4Vc77C8wf4XcdC
SaXmhFW8/TFkEqxsQ4zoTKuN0KjZoq8cj0eeKUaNsvm01wyApP8LU7EK2fWcWckQ2jVdVIkhsjfo
OYFMehsdgPD9J/bSfbcPJNEzTjH9eafkL19x2uWWOZNk1sCxPbUaFk3h5G+na3Yg2Tnuk/3s6Bo3
8Pji/NE36G0vaWdp/IBYe0XzJLFzhijJU422E4c/oSznB7fO/kcZgQhgKoLpH2WqspRO50CAofCk
I6LdKM22tWmjFSmS6/GGWdnPPm4x+qOHKeADMzzPIYh9AgWqnKryMIPqZxmYg9uGgzCCGJU+0Qzq
qtfotV/wGqoi/qKFQNd9hTLmEuv6/dn4a6mvU2lDR+flSYpWEndrjNWUL/eUD+bPbYPuJp9wXNZc
1EU85OaZB4eoXZcYs97IaJFZwQbw1g52yG7qoX8LOT/ixwIWUTkDmzdVywDdo0v1+P/9jObnufh2
7ZkSYlJxM+QEdU2rkUHEPSJAmR82PuNl5idVTgmyHOS9jqIrwOVxjQjwsuS7ec3uskV0D2JMujHt
BpLh++ci3rNfUXxPvHi9lMS8qBzNKlQ+AcwWKT8s9aSL59euN5xGD1gOzWAYgTuc8IAOAB6joImi
wF1rMtIRYCKdyjHe4ZELR1Ch/1/BeetmTk+vBY+dRKxDSgIur9dX1vZU9BKMv3MKX9MTpYDioAsC
gTrUohz4ZJfNVqVcv5Ipqdw4a0szpFVLpINO4/bkahMPgZp/jqSwEpytudtFXrDjuDElBtnVjLCY
j89jyW7bJmsTErISGiJCUaizQebgO1tjTD4OvF67mXzXc/zLubF+Pqedaqbk+E0XObu4n6alzOal
pA3nGT0mKrA9bmWlH9G6Z6A4V+DLR28OAzdYHf6EAWSiCjMgflZbi1D0JGCpQbQ08UnNViMQqin7
TuAfKeXjwVgi/c+ORtVtbUyDl8xI9o/PgO6YPdwOzKszvGKucRzg44IhQxVmIH9TlmZq6ECsh/Wi
JIhx3ol//qwqK6jySIcJgKIAQAhSAGsYYoeAXB6A8mVg7ni91PaqMaxODkTkoM3XUzEhJmxSHPKq
YvuOMDKUbF0y0GY3jAj3VFTXXH+P0Ja4/VHwjUoXrL7D64n4YalWDiaetVLld22rY4gujph8M+3x
g8+UeAjVcVYitSldEfaIt2ext94IjcYY7mnCHEl+JQgpNAwsMkAwHDvf/O5KYDvog+U8H8dVj7KI
MhXDqfr+vqkdrM6NuqsbrtW6JOHH7QzIm33JddTR2gIYgoNalDM5uXyLGrsaQw0R6mlmk4bWzdXX
L572MrNRbifsWPG16IvRzNgN0r0QOfZLlYFG4BKmXnH5D8ud0kxOKHRwi1tblaZ8wqfUKiycCpTA
0Bmi6U4jiY/ZeOCtKXHoFPiJByi3CDhUitYF78JuSXvPYwEv+vSVAsaCGLBs24I9Rb8YVyE4jQEb
JHRGKuF4ibB73mW3hDt84MQ/MV5LpQXp6r5VkQ670qUqrmtCAUH/Y6SOTmCF9myklDRHxsLof9nM
vD+auZmT7q9xf//991PQhBmT8nBw+SOCsvj4kZlnnSjd/X3nR5K6EGHEbro2iwMMbQynUUiblNGF
F3N6ZpjJlLE7KxtvnKixxbPmKhfo6YeJyJcQiWuY00R9hFA4grQ9YbNOVN3YVsWv/DTHxhfDZ8Dx
79uF6070plern6qVzcpSvLn6KJHWKM+Ip734y4/ghmvayEwqMYRiM2r+jRPAag/OmhAycg799KS2
06/5WswfcO6Z4b/0obpBF0foWiEpqj5hoXQksBuMmVxFUjOD+JcTrBSWn2UrQQclFsb7d7pNZfcz
HRbeB9hmmTgmE1PO731AABGo1F5j+2DoouoTaJslPbHNeJ7IUSMuE4lFSHFET6sUNUtv3ty/jZjm
N5SkembtJn3gvWUN9wxV6mobvdmdUnY9dXD414XCGD0pFi9Ri5Elgf1MWGrICXGxjqim37PWOMn7
R0AdXg/QTjpTutGXlXGiD84+lk75k1ZudtjLM1StJwhj9HLSbbExdBIURSBHw8/NpCMRmxuKtxCe
Jxhy7ECKRjILlEP8LCHNDt/ueKChzZpWa2n4VnDCe1oEMsZm44KokgGZNT+237HzbSoVhBbeHcoE
wfssDY3qIAD5Kl635ojW9wFRNeZsO1CzEEc1TwV7E6FF3Cl/gjTIHl1u0f1Q9EgnH9NPSn0Chh4E
Adiw5Yw5YDGz8bZUr2PmUargmZ1WTyJDBkwDuv6aZdn4apcs6D3HDASzWhGyEisW1f5HqVbXZR4o
osUsNIjGOVC3DOyget+i/yQgcJOk1pjXa861LwsBHXaNW2RDUcPKQk8ZLY3sg6yBlv1EbVLmDVN5
grfxPuXOfng7giHSk5Hvf7K1qUodFTLH1GqFBBf30JrbO3o9Ff2ZMmF1z3GEIV2I5DvHUX2I7Tmv
SKzhLNtJZT0yKPjUj6sfGu9EaLcks3AlLAOS7fMW6PMUjvgXsUPGg4rnQ25PuC7+uZv4B3xxtycP
InJtZ7GZXoSOAnPTza6zEuzYanB5SgQXLByn1QV4U3W00F9xmHUE5siULf/KUMXgizjACRdEHrSX
H6AaSaQKGuJwOPbfeopBNln7YKB+D5jZlnc4EphXD0E47dIyu21Qa96LVRa33xnYzmzk66t+NR3t
st66vl9QQcuytA2xkjk7UmkIpRK8aeFMC8DAlp60XcOtXgZR167rMbxjUheHlAAvQmJ9M3MglK8B
bE10Pmcmm0xpEHnYyb5ywqK9q0tfK8fqlautjD1k4Ib+ExgdL7ZexgSbB4Bhc2kutm54gMhlj9zU
xqdhqqVH974DP/ZzjWv2YValRpHxkqJzIdYwtv5A/l3j7UCaOOl39LIm8QIBcKouhG+f7lrFVCpB
+DsU0FGyJg95+p8a8KKP8nh6Jp1qvCCj2NE3KsYowBZMt5y7snveWcKvLTSu6UsBTvBpkKHYHL9u
OHApr3wMnTx/992fGL3lq9p3MLiN181V0YJwsqGTQiwnnl4Q4z13jEvdlMaoapKKiKbHLygHy/7G
pezhs3F+2GHt+eHnaR2qFSGN6QqvEg/eaL5ymsz2LqueoTPZMRqXOWLIQgge5Debtpa05NaYbGCh
2XufdO2tTTvV283auwnC3e/P3Wouo7ekCa9qUffkKGFOsEW/I4cgV2OPVRfmWo31vxcaaD2m7xU7
YLG3n72fXZvaymFi4nl7pUOn+xtp8UDyrFW+ReayWaQ+SXnnMdgfwd4soXBYUSkHTfYLZ4Vo4JL9
bwovWnu3TjBwJGoArywlpaj1XFntuaBR472Y1OFA44+IeTcbRp5yKKBe8CM+XF0zOD6XZcuxP7rB
Eih62Jd2phASxqiZlicNXiZAWWu14cLOnV75Ykyz+wT9C35FJtxgGrmDlULr5zNWUMcCB2mE9uHq
inAoQq/yonaKoSDxBvumTiS1d0T7uWMzxXdZ+vsmzFHLa4U1FIA1yIXFY87J0xLqKyZ+oDfqlfIW
JmcEm8yay1zXM4ycVXExnyksYPBvIA82r2d9NK5Y8A6oS1xNPv5+klxUBEK9LlTl0/ltqSQpySqi
SSX2acMjCwuLHsYzSWX6aqHUrJRSSosVq3ioPnlk6X9Fx0mxm7P38ItVUPmqIEuJUiTT1SZxdQsG
tH+4X+fbn2RhZu4KqDCXX2vZv5iuCx53yofafrv/KKcAzBTg0wi9xbi9E5iq/ks8X6Lqn10F3ie9
CHVmtbUU15DxuvXmThnJbh3qc+A8OcNKWe0EFyXUSQb6uMfPUDH5AjPB4+caERp2R3uDhVpFfSeJ
V0nSUTeUHm2Eqitw8bSjTeVj0ee5P5PEFsH7DldfGzuWo09OXNoTpanpCr9MOGF2Wi60YGB5An2q
EXF0GrEF6jxao27kcaiNInTZjwYZ0pgdaq/g0VEuhd6M9RMaKK/4eCB9Ds208JAY2nMQ+Eq7eIUr
7ldvAVWFs/5qPOrVSLRZ2DcooSChFZ1qM6somQ6fSdogI+sWMlFlbcph61Twgsv2WOIc0QBCG3Yf
WLe2o1QfXyXpqFwMBUExPYH59rRz+N9Pbso6MmSlfMO2QVKq6xG03PJLcH+G/Y7Z4tpHxQqjAD2O
0/ngP1gv+kAg7+ssR6oRLg6TaXmnMOMc01xiZsHlOKpCGLnhQ7tsrKBb+y+cu6gH0j1jqMfgdONt
dtEfPO6xQmR24DLQ90HWUWNw4sC4cCxCxLchZgPoHVnb0rUDpeGSm8cqYSeWU9eOJmH9q2la2YO4
Zf3vXxiD6tmv7QLtOjzzJKzMQcBjeS/fnGv09yUTFCFkENnDlsDFdOJbqNcKCaDVGSnaaPL3Okl0
Nxb6A/YSa711dKPZnFUYn4LT9PyaReZP0gy4dBgmo1xu6sIaI7X1BaAeE5KRgRBqkA7Kty2K8ocY
xkgQvGbHRMgv6n6yKuFkGmmAUX4zsDDxwchmyT2HfVqpE+DQDg4MV4IUH8SHghSze3IRGFlBcJYU
kufv6w8dSrUmRq13NWveOEVaTIRN2JsTQFD3BvW99ACMMDXJnIvBo2MZzGqqhER99+5zAKMkW2yf
uBSvW4tEw1yWCXP6ak9IgO9rkpHMmdky21SHgvyK8ywz8I/9xrBJ+Qad8XruxlXkjc7KLcyfrV/x
Ncf7gP7uAI64B6GhjJaj+vYA9SSZh9l6NvbLVmgB5v9oVS82Vtu1WUq+rVVfe3JxEu5tmSpJCQdW
4fROrePARHmMow/BrPP6vUahV2081Fa6FC8begMrI+02WuqPBUn/AScflR1sw7vTNZscWCR+BqP+
9h5L6cGVsVf+VYdM+Z+FMFzXyKo4Assrft43hP0ijSFH19fNLalHAp/dkRECQhbW62aBt056C+a9
MUysf+vOUfmfR6aIRo4skl22V7NxZahexZu8eu9+Ovi4iiwXFW87kA084Xa/Rsd/w8JPEJSYO7Ma
AMzjOLBElIDbes3iKTgleAmwjSsNhYYGl8vvRsgw2qFZ/u07cXwT+41pb4/p8v9CIO5hoSsVzj2Z
6sEbVladeluUJwrhVK5EX0UCZjiaM0+giQ2kDKD4SYVxb8iWCWgoYR8t6yUSewbnWGRU8fzZrfCP
RGwxzWzDK7eXDLZ5PF+CN8dlu57z7+cCGc6ibPs62bzI8ne99K/CS1o6/E0/3Vvw/e7ia44Zh/2A
MP/KceyllauGAqzdCR5TQp40S3SArQ5eNSjkjx6jDqXzRyw0lpq5P7EFJLwlwUlaHdqO2gYv6ax9
FYc1grX9+k6ZNCK5uk76luJirOjOJyRRv5bDt8e+PMGhws13ZLOw41Yne6vqT9qei+TOxcC9O12U
/omIQwUkLc2UMQAww3VKmD2PGA6TTIqyOXMvYWYPmNArPiKKibf9uremzF0sonlf/AE3uFazdjGe
bFXCf5StsQp6pFUJzT7qpq4qsnZYXf9Po85YCfQ5r50G/dy/g6IVf7NSfbKqMGVssCRq1JL6IYMl
nlxq7UHuI8fvJDocXpnoaSKGqGlPSLGCs13uj2c/mFxAdmxuUGPCvnkhujUVTK7FK/2Mp5UHw5GX
X5lqqIRauaw8YpwGNwAmOu6+CojAUP2SJsGpDU8BgXtGeVm/+ahQLDaLL1uiaKosLuKWNuPKliKO
iFzWL0ENdZAObF7SK4i39DdhocLXajL9Vnm8nInXk9bKzHRhEtx9FepBWxvEJ9ZTEpVpqVMGLcUX
6fnOK9mtHDiZzk1OVUKzlto6iPK6LzA6WHLi+J4D6EoNXcKMnxSMs7FOPgZFnbjtVvqKprBEl2Kn
lQZgRDfHuWZZKPE9WEvRKx9rjgsgLeW1tb/GdTGAnVuSa6aXKDqb8R3G3VoGE6LsTpEb6TuE482k
+gdf96hnnS1Rjb9rzr7MBRqvMw/RQQTKHI4i39fP0fLfGnbZYOPVv0nUhaosFDWAqG7Pv+TxOxKp
W6OE/S0hd06DsoK9vJA8uW181oHQYpRF8cloI+EpwYvQr1egw/hOg4ZgDmbNTCv6yA+pdZV8ZMPl
rkCTxJntf7I2JMeudf2V5O8qNqlPc7rhOLTFIiXsrP07UWbCcjESVkSYyERL6KOci0RJZrs/sNW8
e76r09VrhAyD7c1DEnnwhtFesNSYZx7chThj7cBXsqbGHXDI4xuZ3DU9rWJ/mVvl7nHXR7gyqThn
ugmJxXCR8xL+VTnK0WVkSzuaEkTZmhY4hzjAG7usJ6cfspBMXiTrpGin9wXo2uXGsVO/0hqD3zkC
0Bsjw8PC6FbvIo4m6ngcVA+Cr7lrpMJCA5ezwDBq5PlzGKzfI21iGVM+8QiPPOGSIJjybXhXlfT9
ES2fq8NPjAqNAFJBmPD29nZ3an0vWplWi0mVMcIgn4+4fnqbATOhXDl1FprJJnDadaq3W6Y76PnG
CtWz1TLOvDmJDibwXKNAC+sNXq8KDTD7/iQGjp+8uOe6O5MPP40yS94OTUZ/32EhysQ/Rhqnfu+u
AKXAGBACGb723KXL2aNTVXh4bL8nBuMhhqQgkcSuEtQOjaXQ0QHJWEIf0/DWTkDElqGxRFaGa2b+
uro7E2beCIERozETvvw6IsIs9/FbdDhZYa9E+VIkQYtawg0SnfOSowPofDjSbT0MijQglkLLin40
/JXiwISsNJzVFgJ+qzACw7R/68YLzozAFedqEnPS1FFEpl4Qa27T7oQeyW7bagm2zhm1oWwlCcTG
Ak3PLxF8Nj1MG4BmicW/tUWRa+yvP2OM1B2pbyqMANpoLgeMkTN5Kjk2rJ0kvQoeOxXw6GVmnaBA
EX/m37BEVKdSl5mNUcjLu+Wpdfig54WddjOIQRs8fH0q3mWFy6eTluDkhrNLlghvH22yBFMspXGo
l8lNNirKkTm2MvisVpQnYWnS69C8J4kxxQkjlr9iZ5sB5jgAhij4NkzHCBMPGdBNkMKhR4p4y0h8
5pQs2WChaftXtv5A4GWwp7aZK7OrF1TfcPZZl936vzmKAlWRvlG5Qu5ASdDEAMCnAUMs0t5LPgsc
NMws+ljkxchtnGjunabIjMssxT+u2T54QWpKfrArq4UI5MpPN/YzProNJEgU1RBfzxU5GKemPWBU
OF+rbZT8naL8fbY8ASD1z37Szqq8q/XWWv/hThuBa7OvkkthobxV8BNiOHqlqE5WQkTRkgt9ZWNh
1GNP+7laMTv6rZJh0EhvN5Dk44wTVtSAVpGesUyQ7+JZt19BDhIWAw50cbBOIt+q/uKT6aPLW5zi
7usBS/3pviWNSqfHEgnw08o0TdgqvRn/FAE2PjZvR0Fj5eRhd/al75whFlbT3ztxnkwVn9ENzraY
eroWCvfkc572G3fgHwYXWvHwd7Y9EAwm0U0Rmr4gKdcyA9tP3iyihvICky/JUja5YuvcYr3Il1P6
D7yghe2b0sP60DNN5hhlahdh5QXBYlZcJRTaaXgDGphhf2Ezqio3aOgfb2ViItbxX0gejvdwu80p
4bXfbCupSM+2pglDJPElPnxNbDBzgPgno4pGhw/F9zjkmCBu5l53dcgknW6E05vEL8ofO2uVwQqO
PTJN+ETtq7CYNCUPg5WWgRO6be3+8oOZtRXyNxxBYxjDhnhGP4QDEEBnvOukBk5e9ns1Vackq9nG
Ze1OU/Uje+2pRadmoEIGW6tz6Mw9UNR2fC6pRQD9ytUKyb3SW33FViaSKJQYEDDU0y2zDr3+HTpU
GiQ1tlVzOTk2m9elqep9LXvxNOTfbIda2A67iDoRJnaT7QumLsUCh1X9m9kg0qAFIdTwM+fLOLR2
nVxR+Bk6yTmcB7UmgnCe3xRjTXkKRN9TuX1AmjBFsIWe1WTt//I8oeMB0YZpaQwat/qDQiCPvvZx
EqqkGqwimN5cb/R5CHBXMQpws8plxq2qJeulxcgbEtLheXIgpnPhLj80qUmlhvaE00x3goO9y/bi
gN1GWgUYEJR6aJk188Y4Nyxv4TRRn/UXkK06YQcgdWor35AWFJt1LSd+vHDjJv6xeFo5i+2RNt0f
e7SQy9yLJV/XT2l5yhhzmRlQqV2sVhiIhyDKYvXaf+BvbskOyesskHqG2Su3oyqZzeKtPVKuhpmM
EvUreBd9YsbtQJuVMpAGA1YT6vcGD6dyRS+QDYgF0XI5FKtFhJQtYmx64ChvlOHvyU5BocWZcfgG
eM9jQYvlqCM3Kei/6wnYk1bJLVbfTfXqldTt9Ron5DapU++yZRQUkl0iGxz7R7aGHIeLf17wGvfn
biofYxaARIcVMG1hdLfb4n5LR32fdGZAYabmcrBaMM6os4ttF5prDsNicvRZ097u35Tyjv15gGZ/
DuycIilIB4Sk0LlxVGv7JskCNG5kVEepzejZ5fZHQ1nDBDrt2KV6qqaKgzH5R4Nm03ZfSFYpSGEd
lTtDvLZ7dJYwyhp4smt//gY10nxFeAI0EfScV3B1tIb6+QTNChfR+lujdkmVj9uHGQeCjwnfRJiA
WvIbVBgu9UHpYWJery3CqrEZK1hwOwMsRdvZhT7HnHMjtH8ZlpT1tyTuBf7S0tF8BHUGUM1B7MFd
s4P6lQoqoVcX/wtQLevLXNvhZveNyidedsGvnTg2Gw76IsHvudPVXXuSNrj/+EfD63RQUDRuaRQs
k76bLfLmHl90ez5OTq40/eW69k4jKqNv3hBXh17hPtdWqVlyqD5hZI2zIQojclD14LqrVnC5yKvR
60cdlp3rMGx67Nvdcm+pSOXy0eM2lP5Uu1R1wdV2Puxm1ldsrOFQyA0OMwFFTNsXsSjeQpGuvrce
tn6hAg7VKNQKa+ynXq+PIsHAgIymC/XR01Af586H61gbdVjk7CilxmwhLbU/fdVurxQ1Kq0DCxNF
HLjItJUmw9vvekaz3+DHruBviwGdN4UjaHDdHJJSjleKdVpb42wdVcw6uj4SvSo0I9/W/SVMxeKN
S83MIYmR44sgjacxMnht6qXELHmjAWU+SOJAFDz5dOcdvGIo+clQ5jkqtDrccK/0L7D/3zfTHnA+
ctNk8SHRlKRDiQ/mK1VE9oYMzJZygRcKSV1Ddy7ZeWbq9t3sSJHXEf1p/gsrA5QYuQPBM3rIY8f/
aiZAL48YGblckWWHEInMXr//yJj0E29XC8HgraWLkb+MRg/Wm0TGjSuQzEqqSYc8o9SIZUz7zad9
gd5LUGmjxvKUXjqGWiDPtoWzwptxE6Fyq86hxzV5EixRKGxhEyNo3qLo1/zLw9uVVqLxV0B6sAom
rO2Of7KGKyKt84xzr9NXIpr5k/cb9lZQYY9W1x2oyI7doOiTTKfM2B0OlBPAJ/wdMNYpzpjeJAk8
dQ/jsB5+W1+jXtOn+uOJMnpTtMC1a2uY3WWujobHdEN9JD5V/zZ6wSmR8VEVmK+rlELRBfYy0Z3F
YVN6rtLMbzE7bUiCoEzkaU/HZNsTIjy39cp7lst+R/KWPNSEv8bC3o5QYama/DoLuTVS9oO2FMXX
KVQc8F7QQREQuroJLT4SwI/7twBkRC6LzL50cayW+isV9xPE3pnw8vtV0cg1I+vwP1OzgtT53Zo3
HIWx+pcMfoi4yJVOB69HAVHjDri1s/A9irqy06+u4WETWXa1LfGzc4fQnFizFfgyDBpltJOKCz+8
EL3QF9t1xxBTBLyj8LXo9O4q3KGR9j5POLBUlxVzrvBUljIsU8tpn+iBIWqXt07rZ3cXlL/MvucY
mFNWM7uem3hcqYHn6GtJIuSxNLBx+qBrNn+8GlPY2BZfiXo+Dj8EQmtSoPmbN7q06SR1YqYYO2Xi
Frn+q1P/cF5ecyXZ6DbbhI8UXvp0fgFnN2Mc4M0q220vDSYgPYwGK56EmO/87LJux1a+IatFkVod
/xJtWJhvWwKGHAKFxOk2K5NrdMZREZcoTKTemKHLnHLT+Udc7CVKGkmC8nR++N0+Mk8LTurk+r9f
jee8n4HVON/SIOn4rhYz3m4UVvNPxuOWDUndkW6DWXwZFqcitQqhqUg56H/Le0e7vyOzDpETDDlm
LufQrtLtfe5JTbiHK+2NNoMjitY7iO6GS26KZLtEWc1jTxZLdmSqL/8ZIpNpqCWwPrpb1sBrWwIF
hw39PN4k6T1+oIf2OoA25Fys0H1NHTncDs8Dm+F4yXFPVAG/5ePJaEZsZUWAfRZk2Jm0y5zqLDap
yJI1nkHRm8WeiO1L8ilT/L70k8fMhpS4talXphHevNWUWW/XPMiWPmrGJM76KI0vvfbjKFK/Dpec
AirwO5kjyhaeuVtWrS7xy84lCzjH1DkouCmVaFCg7g3JmfX+3bvZ9oCIoaUJMuhUEChn2MezlTIS
0eCMwqqD+PvCOLulkuUyIlBc8yCdNYm+Q7NJd+vJV8dMVBB+ZmalxTwos/hjmLLZIMaeAZfBcwm+
hVYGzC+0SfgRhGwo5v72MRfMAGmOA29L/PG4wYczN6FwkXfQQfOvkMD9d3MME+tYyAKgT/6XkOZu
YwXU/zgVP5GXlu4RrKhKMnS8IypMVKbAHK7lKhFWiBP7x0RNVI+ylwoHxgfEpaOIvxIdAir0F0qb
XAelunWq0Z9xLDrSBXeN16HdOW9sWtKYTjCe4YszFPG+gPOtPknkBGLXUQ6f9gQ7m0gJUzc2VKWu
TVamS3VMhjRxyhYdwF8fST8yb34dXfoekzO7I8ObQNThL/7AQdTHfe/rqFEbwlVjQSCe2/j8Hekg
oOKr2CEwidwh1OT88Hsqrfb0jNWbqELKz11WCDTfyZ3BXDJWZXefmbn99YfQdU6qIPw9KQvBSRzH
SY/UOb1RmAdk7P2ikeNO6q6ZhIiMszrYeHfqOGv53EoZ1YUvtz/8na14Ws0Mni3SSkoVp/rGMpIL
c/wx4SgxqUWqDUekIU9s6Uezg17/LvnlinCYf8W50O5OlYhucJuT4xAewbLqID7XIup9Z8wSKfnN
JSTSZl9CKX2lBKmN4f/SfP9tJhgvRBch+jj/vEEf/gX5K9Ozp1TleJlvfPvLM7xwMuDX6+a0s2G1
I7KHd67N1XbZWe6ybA9321ol4vcdib17p5VKhoCAx2YGZY3CvfplupzA3PszinB/hH/74MfNDLjm
Y8AI3ak65qjd/1cDAkbMwsjar0HV+WvL6U38YBOJVWTNmk2+PN60QjKbDiIIjWyQ2j9kjWU13R3U
EbfzrDT9xM0oUh15bH7aQzD1cl2Dx4ys54x9S4WwpvQREJbrtD50/yxt+rgeSI8/izUxiQG/GDUn
z/K0JgMUW5AV3GoiEeIHiuXgphUTAMiQA13RIwvyj8aTujj3/HhL/gxp21xf0QtrVidhWb+2vLlB
HJoz3pYWs1nt2HQg9TcgjzLq5q2c+1fVC7HcRrEDK/IoQPGlOvDTuyNG5LwVqrkyX0g3oehPeRtL
M33KkOL2jcPSWHxw47LqgFsKMV0LbChHY+4r9CNfWbre1tXOAeRKG4PFWlEGFKPHSSJOLRXvnorx
ocp0HYUti3gJIqI/8FJpuS2FQ88Mbzknj4Pnf/eQkAiucP9pxLwt2QSPvN8W7g245/40sDW+JhCD
/6iarjLva7CL7+nZUKI1C9Q9HeuixZALI/SdvRe+56opQL7xy//mhyypDFnGMKItWt+NOdXROzaE
J9Pd4VW4hp4Y/kI3gMifvYtHMsJh6JFfmh4EaVPsJr41KSJXuCSEyhRT4JrE8OQ468jzhch9zmKz
B40Ent9G/uSKviLkJAHFllCa1RJi/MhO0NhsqeqYoj/iVb7tqXInyi0uMhsS5oFpMq0bIJMBoyos
Lmy2s9Rg6VOopbpHeq8H1+hDSygmrN8tURoTr+ns26xm0sMv732T/XWtojTOMmBCk+eL5hBpQDaI
bTyPpdsHc+BQLsI4epK1JOcpo4sCVWZPF/z/O9HsoSwYMHK78zRtjoQgR9v8sCp+yBAPA4P8wpSj
zgaidWaEjNOihmWE3PHAI6Whx/xdmjkaCWx8jD0mDLJCKKjjVffWpG15ZJZ8nCSvYDyE4kNnNI2R
yTgdpa0XEdI7qZcOaGZaySYTxeaI6QYkwGsOyiQJv/lYkJQjIVfNHcjG7GCa2sUpWvYM2cK8aJda
NfWtShSgEgtErgFbV8MlHk2zsy5hxIA8lNXntO/kkbRj0eViSFSXwGWzOLnc2DfYbOKURjhTbzfk
VkXAkqh8CaZbUREU0ch7M25g4jhHaPvmhoN308LiaP6j8f6PmUO5moQ2jFb01cjkDHOzYS8tuLs9
9UorKRFBE5QvHquHgp/aQz9NdHfud2zf6Hd5AEpSf8yAONuiXgIcQSNauRK+d6hOazoxuIU7c45N
qa4d+v/6QgCKGj5/BsCD+acdH6PXJNPBif0Tsb/4I0aDUhgm3Mi2qVuXoX9eAdOw11Ed/NZ3jWrU
2+FW8qbEjZemPBNyX6auxMrevdzfwG9BlDZKDJLtcfmkau6y1HvKG1XaiItTHDjQ4mAFgTJLyuiz
GRpOgA7NhQjRH0H63OIVTyYWLwypyG0VlfTmPc07/e88vf3LLNkB76I0PZa6SJJCYOa00R4uw30C
17cS1D6FIv85MnGcDzC1K8H6KMPTPYoHONqTTmi0evGa/gT0X1ppGxTYWtBo3FQ71jqmGsC+3Z8Z
yu7Nl7putrJw2jRZUTL+v3QGIyiPNDIYwWbRvgjzRwJ7pIrqOC0T+o5GagJE4sS5KKh076+uwQG7
eXy7+5FGKyA1rPSDdvqHk+fn8xaEC+JjFZ6CoHib68/HeBO/hniU1dBhwo8rTxphG5RDmUYOqXCr
DJH59m5PTJCGQoKF1iLBQlY2cdaAPgl/udmJDwEbFCymHM/Z1gZy3IRbd9Xn4vYvpj/dSnleyPo3
oEVNfDi5gaGnApsUmgj0VzkRjr1TLFLU17l78fEOGk3l9ulB4L5egAfYBXNcqctFQU5dmEJal45J
YOmD4TGDtBUgapERuiULQ2hEPxXU7pp9XMsgt5zKswPK+ZZ1N4YztNQI1sos71ae/Jlbn8rRiwq/
15b1+kto1qZ05MrTKw9kYVwJn8q3BA22Pt4CpoH7cn2bgI9s9PNx7NCbHMK1Zc6dUSTPyQFNmT9F
MvgdfY/qVknAm80LyG9Iyv+qxbQNsL0dFavphBYlILgIte2q7FUus6yv1rI0yMNFhNxsPEw4Rd4R
ufyvM8KvZo4Dbba6afUonAZS0bXhYIagCV9ywzTEeRG8cuhr7jmN1uMOdTTi+yOC+YmkkcVcIMSO
hXpetMKrMVJiA6U2cU5GXgRfirSyYuJfnbqFQZOeODBeN8+H8uP314YX2tN/kWu7mL3HPmiunXCR
CM2U4oxzN0gjZgilesOP1m26Y3yXk+rq+neMwoSoP2rZbdpPIAOPn88jQB9XyPqKKfgINxDrm5ik
8oof44L7ESvvfkjOJDN+87tGw8aKp6UvltzkgzeKFOG68ZOR62bJ464Kj9n3DDZk6FEMYO3aBpRQ
7tdChPWw49MkxzvcCAyEpRdhF2LTFucepCz4JGMbakWAtpIS/TIC5zdu6ak4a+ze0kJcZCTkHYFd
bN/C4//Z0321U9F4kvWDbmoXNJvWyDNByK6M2TBoGE9TAZ7q4w82DVY+TQtNzg1hY22JAk3VgkuH
xWTGgzu97M4SJ5aal7ee4pzituchFyofyjk0OYxggXpjY0xY+ckRkGHwKYxg67kTPNWZGlsrEzXb
5Y3kzGJUFDXA6UvbYxeJjuqvAyEOlg7iot8QMd6Ubtd6/ZTgbtB0240O86WuJeF9BvYQxmnQDgRP
kF9E2mE9SpTDyQchZp/kWPk77wRRO5mCGf2IrVuGPDXTuWEKLHgD0mi/HmPj6Fu3i9xiJItqO4Wg
yauCn1de636npPoAuRwao3QvFT9B74rDfAipmWhg/1cVlvObh+Bb6JwzsCH2hBTGIUJUbFiWES06
aE7YBPhWKuVORcNMHr2LZqYNMg/VCFEBLZkrf8imsfDb1nTOkYHCe1yTJXLYksTr7KyRR8vDaYIv
o30c6SsKT/A1ccMDMbOKsgBTlksh6N5JUoMzebP2cfdA/60JYdL1HkveElA9n12qQfQcWQFOBfhf
EvylzwC4GLnpnmuULHqdswCxIPGMXyFQ6F2zASNiSUKPv/a7kbz+0HRTJYq9IWEpwzWW/0pJiUv1
J2bdY+jVZ6gP4vbftbbp/YmMSHl1/8Hvwl8DVqGdgVVr2/uN7HFs93+kykUhN5a1apJGf0mqu/ue
nW84ffllra3C7UaqNMrO5/Hmypl6ehS5QUuB0On49SzXQebx81wUBJ0dKE9WA1+60gzCHuBloKMN
TRIS36n3PMhHsExm7t17a6KDBChrkKR3fujQDPDWPyeCSJ85Qch4ewfECU9PymloX8sM0nuFl2KQ
kJf2d3uMCdzg0xsRSVqz+j0kBDybeqCjeU/mUdMU0SrNHNuKsFSNbjYlryiL8V8WR4dnOeHajR6u
L6v8BY5FbE7QZql8pMUuxlkyZonjmGZ+lOoVDusGckUC2Jm0ynGFXlGSPzRcIWxKRNnJERhBRFfI
Cf8iTIvwJIdO5pG2Bf3HEXg9a1ZbRXLDoZjBLGAGoL/Oj8nfd8YbCl2bSdyDBR5Zy6Io5WOOWsmU
L7S3eh81m8twV8AuyFn/PrTVWciQbM+fYiDqXjkf0Os9Jdmy7/IACL2H1xoCQaEOF78IAuNplxk8
G/M8m7kRkHKBlXNKgabBfwaUoUVHN0t6MnzW/7+4GOSzWUuBz0BV59cNH8cghjrfPSYBLpFa6+R4
3UDXIgGnrYQeq/N4L0ujWyRlmTRSMOYiGol3mlf6bdZgtuSjcxpVzf6j/mToW5TiJ8xE68dAsqmr
EEhqr7+7dTgmS1QcptaA/qM2+2iE8K4O0i980+sO4yF6sfTWO/s8yhoPpfBWLfUQieQVjUI7qbX3
km8opn1kTY/16twaOD3A4UzFqoIYzXNFJsOkokEzbhHkgunULy6aDVSuAXWPriaYBp14lJG1t9jb
0ED6c8gGpL+b/oZW8v8u7eI7CAItJozZFy/TXlLvB0NYRlFVwHjdje64D7VHi1slyXr3DQFZFxoE
9DQiFV2/jLP86WQl0pCyp8yy01tLfjFVMBxIaUnxmXej+Ozx3+/DbOTFrJcOLElb4m9iV1rjhrNb
nzCtz45EWJSnEUYqv7Lmpx/c27sQb6u3tVDoTldQlUoPD0RmufAvSB7KEMEedmpUbG5GrVrgexZd
4F63S14r2rG7WGKf/P211eFK6vVWfc9msre/zrZrPXmoajsYN5Atr/8aN1xYQZy1hTIOdfIxCqd9
jOm5r/q0A/rJ1UFMLlI0LNSRclNLEbpeZft6RL1Q3vRhAER/xfYJhgxGHr/7I8a+oVzYQCq0ptXX
UtsnEpPGvwaxFeHywQRjl31aEJ4ggmXoGZAi20wEwv/QUX6gEeNBhz7ejsTyXUc4WdP6EVj2rerb
wddxdhagvk8h/dlaFaiUR3ytu50kYm4AiHoi0g2GXOmNRPR06LrX6vz5NYd+zhPbexoanxfyyy0G
0JGZwJdSv8KFHmxoS9CETsmm/uEdVDqzUuyJrU/wZq03nR+eWz2SvkIY28mOdnCvwBpGLkwgBjRM
Iaeq7hNicyV1QaAaceQKDy35JMfAPg+rmR47kIiTL65QTCt+kpr6PfNCg/ELSc0J867DuCoQIXfh
nVQ6SCte9FNMB1mKmfeJ8yPCbQR51CGjbbtPn9cupMdCnFlnB1EEM2Q2f+x4vCxOBrmGBuaqgar5
0lJ5BT11DCEA01uF5FVz3qG5lRlrkrPs251Yl2GcxMUtxtBF2TPs2TWwqS+F4tbKuE0nIOUAOF1P
XjkYHuamTHi0NNzCEdWPbNm8Rh7maY/x3qnsny78CoFrYQbP7l8V23BE52aQIAV2YkpKaEg3XIjx
0rb72kizEve8Z+zUJ8BRoKrTtCW5uzoZYO2O5LF8sjjv4ebAPAgo+lj58j8ALyMpTuAry42xwdDw
p/Nb4QqmKT/NH0KQt2qoX7usWSx5I0tdHst+pqtCReGqiFowg8ugVxQ5Hn6k3va/4Cw1hUgsl8yh
1x7ne7/V+jz1DVvjxHlChvCw2eSW+dyzBzuXdqYiMuqidANc9QjkJ4+ajsRiyX5/t4NBN+Xzhbch
m9SWgEXSXbrHKTylH5IQZx7fduVedOOEHDThdpjJGnbNjd2kGXYnHDlPJSLSvzgBW/byiEtnizke
03hCrm13jBWjYxUoJeueuRLQkHh7Ofo7JUzriGfQx/XMgIbVczVOoeX0+a689UgWs+6fxvZtpNh9
MR0tFn+owRe37E4eV4tNpb3dLG5LBBWGRvY5zkqJ+cisKw2Bp4mnQd3IqTonl0vf4o6TMVmzilDQ
/UkvCOMr40xWXFoW7nNuJkCH/K2yQIn5wLaj9Z9lmSPBgCQptATm63v2Le541buh7NDxIuSe0VyB
94IM/ou824ruvWXj87H/BoYlbea3Uply77WLtKGPc40PqO5XZouvPWQyKbkExq1t2UgAKVr7QEEF
92RPdWxTcuHNtpSRvKaDYnJ7y9sU/L/ryMIXrsTnYcGXyRKxvvyWEBBCICwOEyTakia5zusAzGay
Y+21Kh5BDZmIqN66BRzyl0JgajhuT6aFRCdXDNcbIDjyjI8DqU4kNNBpaRbryT1BD1KuCq4VTuMP
65dDE0xIuS/K/4hSz+hDK2/XRkODNDbkkNY1pZ6LNFZp367AaJZuFrhgxQPGwV2TWfgKBvqEtRuP
2T5odZT9em+gS6Otc/DafT+Cqkv1cIzbflox90tBq9eNlk4qV9OVWIFHZNfZUw1rJauNBtvb0Flp
bNnujVHlMzskYcgBO7PCJKVbl/74vMxFrYRfLTmpwUwqqCP5ujIr/wPP80Vc+qvaJVwW6cj4Liv5
j0GJ72s1/QFfwI75T6NoezUkMxzAY+wZ/ZAQY4tbInHn41e0FJJjHDvjvr8SM7TL9Tcq/3vcEyyJ
Yh6TTkJ5KR/Tyrt6n5tvGaf1yK4UQ+5IU0PnLNXJbFNAXTVMBTNiuXkliz0gK8lXikKFIHLv8A44
Mde95Q5TP1gVAobzGOI2oeYs3CMlWmy15jG3za+468zmURuUwyzGLBmYTflpSnuBN3oW0wJbysLI
J28MVXaECvA+uT7ZmuPZH1i3c+a5daBU36F4+HT8hPHNUotbbZ1XUh/4w8lGo3vUSdj1RFd/7TGS
MUJGIJXsj2qbPh5/MayjrP0i+TA/ouQ14PcTByp8KsRebCvf1g09oRyMH9FOXjk675dr8UC42hEK
1PwLXgSnAkiWeW9Q3HkFXyyJKx2lUoqNHTpg5aN0HzCQa3OqvouAvLN/NRLAX1nhb84s2qFWSVu4
j14fT7iX/b8UN2MUsGkm+aS1RWUFvkkTzTg3Wkv1A96xAeVCDKl/3BkolMeCKFxZITeFswFu4BIH
1XQ6/pI+XKetdlcdvxz6YtelVwOMxKzMLPPqXH+vc7lg4MluCAFwu0168F6HItlMISp7jB0KtyEC
hWpFcnNtLWLO8Lur4o6h6XkpRGjT0LegEOgM2GNFouI9HtHEZ9NrmFrgRxsyydgst6ra3LwDGYoz
OFLZQ/In+42YjB31zRklDnw6M9DwDzPd/mjyBlm8BSHZHM1dzDaJ4CtCcwn+RbCEv2IZ3h67wXu9
cS47YdBFrT7LBwxy9HDzRxuKyeLIi0NUzlR6YgHqaM7BUy9kNbuaHN4HOK0dxObFgGeAI8taYFNK
vN7NNQPLnmUaFQPMmmw48I7GfIyaOp3ZfuwQ/WxZIWGID1f0u8cKOtPEdso2J91ma3tjR9eqb8aU
tA7OwcLxDqAyC7qRb+xSIWvFjTEewABsQ9f5E2gcg+y1OMJlP3eoLyeOec8KrtUXUfi3bONAXclk
QCMtykUoXsngNWBLmzfDu+4TXGeu94jKAPdmvgstubm3Tln+RMUpR6vN4YbRvgSNAnSfqVDFp3rZ
lQjPFz5zp3AQrvf/HFpoi0osYC7T97iBnWZMRKoVeayH1S1hsnh1E8UCqEYaxdgCH0OOVIMg2Ap+
3AgZNlUuh4VWPnR3JXRR0pOZGKx/mL8zzAlpylm1BWWPEfHMaVPvRC74C19F0MDQ5+B9eNCXouQG
yg/ksZzYm8Uq8oGIaVJg6TrvjqYt0nzvy6Vl6zNukUp8yx0YwpMM1OXtDvJ8r2qLtc3oA1cQAbOF
V9T3vIUJAxDbcp2IMMBbaqkkWPKkclpsnxRjbt4GEV8hK3uROP+my+OLWCl6lsKSH8eEnGqEuODo
1xDqcYoF/G+5M9Ze90vZI/b0Ybx+JQiM6yRk/AewVzae0VHvRvmqvkPhc+wgCpTxQW9NJZ3/HyA0
mnReZ8VJratt8LztcMEgmXV7IDzhfLg5Iord+7cZz/Jcllle5UMnpU/pmexp7/oZDm3E907lGL29
e6gNVY3gW/0dSQmh7Bf45JcNsMjxzKPMevL/K7vmHfAnn1TJEBc7DD3h8gkFLE7MirNBP9BUF/xU
w0+8nbBKCAhZ/5uZiFMZufWHi8QMvHVHHkVLC9e0gtqY+LS8VnkBAxhtnLoLFfGXfB1PvWMzG80p
wDEW2gPz59YZ7EhTLxgxH2xhnsIofi4kwDry42nO4jZDDlTEkarIyTIdfNQW0oLM3YkoDgV5V9ZZ
9w50MAMr9dKRhzs1YiXOYRsI/Rd+FrPxGPmDbOx0ThH5ghsLNXAe7W8NrxmKmba4hem5BGYQrg34
dBPvDO7EzIxMpnn/ZDaUAyFPx+b4mPH3qP7TkTXrGPl7TCImnZpIET1XCVQgdO7JbUalFwr+CzJn
RGiUBj7Yo1MH6OS1O+Zf51WwkDiNBDLDpuqVJFyiE2zC5hgbIU8LNBxx1GGRHSy+JSevsH2RXv1Q
HkErBH0aQTIZssgbPutM2sM3cctr1BXk+PD+q6ThYROB8zn59Xe2HT1F4ZLrxIsPdiJ4IdlZHBcv
N7sNulomDaH6kmW62MJ4suKCMrlvqnavuFRyIguUNifzW7aHfD4pGLhLuD1Zi1Q48Zp0JrKHI1Jf
1HkTLymPEnNrxn3ZU530XzkXZq4sIWAJ+DtSajHvaZhmag77aKEKrM1dJs3LgHfKpUnSfFwYy3JP
xNdhmHtc1rzoQ3do5CQKcq2ByeeU6xnswpAk42B0BDaHyv3Ee8xh+Erc2fH8qwktV8l7lIg4P4Eq
cs8Vu8rDhkVhTxqqiu9Tqfzua0Esysr/Kzi0/RMWc5SVtF2KQIPh8Bklsz83N5gZcsT9vj6psn/F
tkbYBb7yS3chglbjBBS0lmFg3nTt4qpNAXjPa5HarAbVnQYZvjPJ9NrWrrL5RjqYJ9sUvvJjxxxD
y0Wgj0MIY+pkYVFOChsfNqnErNRt6pZbZ2n5I4tTOR5HsHK4ig/j/zIwkMTT5uxrCIZyQ0mZzpet
ne45db2R31Gd+r/dnpVYMabpmmvZ6808XNg7hBW6BUytrSq4qIUHARkK+D1r4h8g24ssl0QuDlp+
ltr9uATSdf+df5ykFzLWipQaJUZSZ+5IVPUDFUp45gf9UpuNSgdru8XuhWrZNLQOP6Q8rZlX4Hle
/UgKlQUYGM/b0b8Seg+opIfll0SnuFXXD6qgNKpT/12fYPKyViKGQFfSBw7T24HSpNxtoNYCahrl
OU0Urx1h/kMaIfe9e+WVVXAbOtvnKw4d0vjieKbyF333x0qQCh7CKDn4cIfi8sF/+5T0f1VBY6ZT
Fbvyy8qyPu8MOxBqYgJuaISnRiqMLd55rFXXVUUg1SwEWVhqOx8joxjkt8JSvATzOyP7VLE+8JiM
KfPjwrm/3bjf+EhGZK07LR1CPnoSBkFOSUnOk2HyZSnTSiQ4yZd+ojjnZ9dgC+HZ4GPwKfv5KHeV
0fc4xoMUzP+x0033ln1TUcU5kn2aOH9yFBx+Rch6PmVLaVVrZ1xxWBDt9tSkaUNUv79DNVb+PMGZ
FkUCB8UHCIMm/dfJRxRgLHxFoeL4NnjZOIAqo3lYk0OCVWyS+tUtm4jvsRi1lpo5SyeNOs3g1Fiq
pNZkoT4LU+80Tjm205XSiUB0NVoh2hZd0ygnKS7hg0Ea6//mhe2NTAEQiErAhwxxZPA35iNys//p
AdtrxhPbsOLYwhaAKKPYAyE8+fx9RT+2Xo7jRn2Mkw0SLZ4KMtFHAZe6opLJbCL7TkjK0bwPs0o0
2RzVY0TMXHuGoUi3Pa8Pi2bFEQt/5I9gJnK1nDe5/CwLYkB/MzapjbnrrMNJo28USxuNC7CbCFkG
U/f3aW1VpYPzMBLtCJv/xT/5iodglvp4yqOhETGgcQucI9fHkDjlFcQ6p1w1KqLK9f2MxwbOWiv2
5o7/htnVS0UdetZHAJ4Eec3l1e1/NYv7cg37Z5TLQs7z8Czy7Jge6bZic20vrgVCsHPneFDUqdOW
Lj1c1CbN2IIglz/PbhSWDA5u6gBXOVV9CkywuU4d3nUZ1CEV6zzWU0cVnHKHr/cE16JmSKlb9ydp
J7FboVhV/0n4xLkCWF6tHFXdULRLBtLxsIXpVqmfIfJUOySh6Hx3U4i33Ez0mgOX+ZOgrUdGNTHt
fUDS4NKo8sTwK609zYtAmhBAfWgb3OCwjazaloavaBSfu09T3H1JmY7eIaWohAzeyIB0zFYOaQEF
DKwbCeVLk47tqbl6aslOrj7NJo4KX1unLSD9XKPyZhnh+PER9vq9tM3zC1nDD0e8gDVEgs+NIAMM
3wzLdGxZTCC7VFodof75cnoKQrUSFyGIEz3VRMY/XyqbKNmIj3c2d5feCsI/vs/FqUgOOtJQVOAf
VySrAwP/aTwqsyJecKmKCHblb/FvP2OZxwpApt7Km+TI3prKSmmh3YA3D+55J3d9+xi1ITF8QrYo
hIIQ4rumSIgd7aQhtW65ReruUR4RSRr/CuBTndS1uczzl0OPZXflWpUQkqYbWqnxxH2XgA7UNa01
NMHaHxlWJwmlJmIr7VqQJV3TaX7++cne4Fo3VtSd3IEx5xeY4IgI/uifWvWC1cFPIkB+6qGTbJT+
BBNGwVJvQTLIQb+/HG1y2FBmiN7hJGKLf9P20ap9KUaE6VrRrTeoZSC9JolxCiZbBYLhpL9KBs2c
D4p95cm1YYH8ryUj1egPWsstz5A5KfmDvh/hQMcJXxFAJ0pMVwiyMBg8mgwhaPEKbQIg3FHkEaTN
wR8s/RYkzU0JIc90xIX+Z5mRsvJWKFdf4izZOOmlEPJIq8YzOEIYR86FcUq1OITl9TwxKlpZGCum
Ob0nLj1ATCNR5VfZMjwU0ueQH4DeWLQRxU+UgIDa3EW5U/l6k95r7fHISxRoggV52irU6smI+UG4
J6Uo6ArDo/h2tBJgYXw0rjw5YjqKaDBdRoA6+WKTU4FErsDmxPo7oeHPWvjESQLABDCPooo68lLq
im9tRn4A89UGwqi61WOK9Wv9gUZjeUdRcqCFInCuojWqp3vWpwaUY64+Y2kNtVtmB+lHMVEU4Uj1
YlG6xoS2dg/+ak+Q0pn+zH5Zi/u0U0xAm0AdajVNEx0HdaS8TNQqa1kTqbX7fGwZJPiE1jLcKEmg
ZQgYtFOp5GAYH8x9UiB9Usz8rbjGFXGpa4LYXYi3d1aHA+WR3Z+I0WXZ/jc5K4bys6mfIJnv8eom
lk0e6TuESW6nTookX74t3fUzEO3LXKqOix4b8Jq4Z5UsjBXZxsT2QiVNU/Zx5BudcGhpZavWCSVX
AWdA0lO7CEcxP3Yff8BO26EYp0s/USY8ikES6ipliJBsI1+0urMOiSXbv8l9+nNk6J13vNep/5r8
PeQeQuehByWCS1Vy2P22tDskqY+7kCmOrYJCU3C1l4QKVEOJsQnPoFpeHp7mqy1+8OEnI7DZUQK2
mn1NBaCe0WwfqXUKG5cmXqi8aCP2krv0G2/wNDDNti0Cmc7t/cf1gfsRhE/LxfMPYSFgc1cYTCu4
Q6IA3M/TUoqJ0YqTzU+rHWO4V1whBWyedL3sUZvM2mnTt1pTGMJIqENpAH3zXZYyJqTHbea882Xb
R+wFLvqluxQxvcoXz8zBVKpCNZBGxvOnx0Gcawoque/nB0PnnhUjUTHZipdE+tbOeS5z3ow3Y9ju
QVKvQGKKfmNsA1Rw8OuCs4bHTl1J4IxHles2yT8tQeEr5NMVA6GXaSdHZ62xXjTe2J1Gg7E6FAQV
hnrKdHTA7zgkiLSY6PhicGSbO/DxbfV2gWf5LyxbvC9Mv1ueO1/MDUVcnhLR0bbaB2UCPBSeM1g3
GImFNcrw6/M0N4lLcEnN6fJvu8boPVOGkOrLt8P2Ds5kRr2UxURUHNYIcuIVmlh0mEy+VBX8dTs/
zYiB6hv9UGquEvR77vM2q3l1HRET99sqxBLpQ/aHMVt9qnN91mwafGUJcbNnlrnhYJqBaSlSqn/I
kgIIJR1oGVFTu7tys5qjxa5Mesx5pSEY/qtAingVFkZUO1OXbTQR7IB1ctNQ7I3/3NINHPRphx10
7mTmqGpiAEuUrFfUpyLToVOjxjYYhfGH0OrW0sWA+9aON0tzBQUNJ9vWyx46m8DxhtXr5lCKP315
OLOoxO/0tADdjNOPi7gWCxFDBO62Ay88v91uf/FKoYCRocqazARu80IhRTOV7bnzt+9oDncD4Awd
oP8BC2dn1xveEXAAyFUAR5qfFdOTFftkQRHhpoND3qdRchHA7okkyWyg7IWbslgjlWVJKePfDSi3
v9TYMrsDUoEqPgdmA6gYamLgmhLaL04jYyNJBkUHA073LHhl3WHP2q3U9hokGQtu0f/O+aqiA6v3
3tWXaB5PR5wsZ8qg/SCcmiyQywb8i0ReX05fpuV9ppUT0vHOSBLntB22Dc4YN5VhKod4q5ejLtQo
9itBymkwaYmB746U+Asl8mTmsTSdR9cluZCuqx68hb/nveZeGDnGsucygkQKOQJ3Z/wZ+UwjSgb5
RTPOtYZr+8ejFUaZQJ7Ph+mnnsBYjlLJoV/f3cpQR37le93Op995BE8CZcUEyP9nnftJqlCgFZbD
qq3hIfMynLXmPEu1r8GPtfIpqwoY6CLm9kSzgJuChnA+iQNRGvjg5JtehMqpnIOcHSeB4fneATRd
ojdLpv2p0LP8mp/NjM17gyKf7QUF5fY7gS3Y9BIlUrhaaN+Vc1jFX3ufVGhFdGs/FD7AZTjWj3MB
e2xFQkEkuNSjbeq1Oa+5xCYVogJjQDVIGth/NwxFCuNYPjSd3GrWEWRdgy+3A2EAODODP+MBUunO
M1aPCYyS9NAt2U8fwhB9ZJaZPAbx2yAJhCePSfYB7RU2/P7APFyefzU9FbgbGRq+uOegaNNfsWym
5dnnQ7Oi5ddRYOvNWx4FJcQKxwsvpOfNk0ZKP5OjkH5qLX2IGjNwV96mieLpN7F1FCWSuMc+14a5
dDvkWBRXD1yiAiffSrl/8ns94nVfFj6IAV+92wXT07/DoEC4l+FpLnFc33eZjSUdDDkUl6qSR6MR
PjETXf7GVRxym5Mc2nFWNEyk6cuikjV6Uvw7EFPYg3HygnHQ3ZYGyqgyYS2AFpqQ6azC/JoBCbXO
JmGu7ooRoY/kacavyf/yLK0o6LL5kVaLZzaw+S8Jmku1lqj7wX2uGkWvIMJQXykXwXFbjdJihIvw
LkKfbYTuVxkDDuvBuA8kJUmz/VBFGc+6JQSNLro7jBOv7KCNL9yNJjme2nck3aCthSPLjEIxXdWS
sCuhQNn9qOQjazMAjzj74LGvlfXlpq8OkDADKS+gtAiAc17IMjFxiNnHgdmUk4bnSk7G9xkTF+Pm
gSRPIzwu4ib8aNCwNvsEJ33LDEvL4Np+n0T4BdfDpmmHS24ZrzN08KKD2Ya1lJBZ/QT7/BJCzIUI
y9uX6nUZtY0fst6G1/i0Rjf8iOK8JtMZ835vubOl7nie2V2MsL0Z8FBUSE42mNF0mDqEjGWkScek
ikpAIfQ5zmMgkTRZ4VdPmJ59Udv81XPGt7zhAo9dMNAW+iNoLtkO/+Pgk0g2b9Cew8+4jHMHcFtW
hTXp10nXv06FrVcsVhpIvXiAD3JcKbiR/J+Ne6eJvKPBo6o8Hg3PqURMWc1WITV4on2a4ylVw4hE
yryMg4voPCY5eNEYXV88dR9Byk/OhA0UdZGUv0a2c5/9bcUFa2b93ZWIe8AFIfLERdYB5lH7HqmW
gjs+7ZepxUUo7nzcx3fWVJACGMQ6cT4Mu7XAAbXXrbVWFsH5F3EILURDcdTTPqppNmVRnM6XxgHq
Z2s+ki5b0cJZOyhEtGkbA1qea+2vkhbAk8Ob4SntbVK3dg/DOw0aDdClhi7Py+8R4m1OuXLgYRMV
0eN8Rd78oXbBj2PjLfChOEDbecLjxRzxqsliaw3wEjiLMVwojgP+ywB6WqdbITSu+TECHejNAVF+
gelBmArC6pen6F4nNlDVr6z+4iuO/QZ8TwVQn8ZnNaC8ZsfAvD+WHvXudmVM+7yLNdsMjuY3p7Bp
ai2Wp6cSPlQ4eIjaEjvoZ2s9e3DmD8uxz+EFrxoz8DYp94uhi3Z8s/L0RFGsKbfYw2xRVbiBe4/d
K4yp4AGnryJjHrXn5mb3XdOpnZoecvW1Z9tA2PUbFHqsGtoQBtCiR2NdbJo1b5NTaHPU+DWihY4a
fZ9y8qglMHZlbfTzAuj9DziVWp0FyohQEikN7O3uvRCll9mtlT0oElz+18xNOJqTeVifCevJibld
QLg4qqhsFn0Hvluffzh4VcJIwWfKFcZunOrlmGs/zoFbMD2SaGcff0bxqUeTXx4w18CEAeGiR980
WjW9luAaD4FJbuHWFnOYLH3eSQKk6ilyQnPJPZVZbbJOdvF95PCpwk7+DphcAg+ot0ff1V1myxui
jW0rYEqQNOuT6PFCxiDs+vmWQm8SZk5IiCvlVfIn97p3xL2NzlprV6KUTcFYd00gBWR24o91JTGu
KwBv2H7R+ykNDDKCfcN+B6ToXRPmQPncRUFYDCXbVA/JLjI56YkSGr5Jni4V5xlz8Td3jyW/BzQ8
ZHZ2593NVV5j07CqS0njxNo2SZlbfFCfsSnCFJvmEG+KVIrrOR03yiU+VnUvjJuVPdEgyJcHQdPl
KEGd9lbUTp1e8wE4BtWBm3OlXM4V/Z6ZkIZKSXixgCaO+A5uzgJSVhZCJviPNqu012MbUqNV64J+
hUm73jhL1XqfX+xelWcj+Xmlx7SY42y8NhWwmNGw9MGs8vKjB9pvTP9X4/rA75lBUwgICZtZ5VBU
W1Zty/GlNysrYn8+2kZjNeSmuLfZCC+cXAn93X9rbUc8WBYImiZHLGJuPjTI1282cEyygYwxi3Jo
tEJ3s89brf7Hbg5qNzKIhlr72GE8fg/A6BX1V9vGaU9YeL3T3qZRvTy14TPJ5lMUKaWNMs1Ye9xV
mypFgrJDYeeV19H11T6WRNWa3TtEucYN242xJRKx60JPcFgVFajUWW219i4ZhNW0Yzc7qe8ojzww
6M/KKuJ1PUfjS3QKYxh50xWA5XK/1gBYUSjxPBSA5qgFhn8ywMS7RP3XbLVLxyZZbMvkH7y+aaNz
T2Fs1wpSHwIAUZi1q8PRzyzlMHEM5Ni2bHuaBFQA0nWujJCWzo1/UxdmXyk8q+yx/0n6z3v4e24a
Vf6K6rjCtkNYceWGbj3lzd5U5OUXzhNdnxqM8TR1Bpoz839HYtm7CUJQo3+k1ANpys/BTYceuXps
i871aL62gz/vzgXIQ+xGvLS/JGINnAe/4W79IWlwItpFMd3H6I4ATkv12qDEeMqhWRXT2riLD6QO
09n60I3nJ4P0FKEZDyrZ5Rk6xExgy/KNGc+QfeSlUl0vUgQt7qtizW/ar0Hywj9vTtS+DtTRYAiv
OU330ihZ7BGakdauptOmkU1NWGLvT0hmmn44UishIlMhpOZug7rk5F8h4magjuvPkH+waUAfZz89
6WusAlNmi0iel9fHHPG8Q0O68lx3/fMlZof5DrvfhzjEgzIRd9MJquyk1c87gjpeclne46YkCMX+
eZMNldk1evfDocuXxBa66k0EbUQ8gUPfBTZkvI4uUyPZLa2XU+xM//tiO7vMndk/m5cdSQ9TwlXr
LwbfyEHS/w2rvA+VgeRmEtoRgvV7O/pCOeRsebh+xh+E21OGZBECLgnhh1g5MybqQ9jIp///FZ84
raI8pPFeZZRRulchR8MGk4FmfS6SRB+KR0ShIdmV8ZjweInn0Ivw/2Klvi5r5oetYdcwK4ABlAMS
Ty7oMxMvycul6yHtx91gwh9GRh/VFiwCTYF1bBpADxI7S6juqtmlg3HcLhct8JyiNyTFjF7yF57+
WTSYfrbhEZZcdJaoQyV4GXlaNXQPrPLn7lBQ0wUEcrwi+PJMgv8aMavoSty/kN92CpRqaV1puU5K
dfnB067PlpZgGpxiFhKDUE4/zD6tIfnxAqdPk7mL10dPIq+XOShOi52knzMTcPGF+7rxqioVJPde
OvUEmxPra6nhv8r8O+hpCaXbmDXLAWgbPY9ns+RZI1SLCrFJCim3ae65rg4UkXMK9WZ8o0QmIxr7
6e+BMZH8PlaQ7dZvSbOGnUE96G/YVyD2GMtCoOKN6SY+BinmvhVdxBlSNWj5RXwj2SjoGnApnMQV
q4P6IiWnxW4dJ2UZwipCrAQCQwWLR9EN2UEKjpuHBALpQd18I+IY8ZMAGe97dLwwTlEmjfoqimy9
Q/A3PgZzLfk9J6ezCRRNtK6e3V9mPQVcW6vcvwFhayMSfpSzYd5JALd74jYYDJ7hCUAC60WYuMfY
uusX7r+vQ/YqeK/tEcjAzJsOlPu+ai5Uz8VSOykmguA36W9/t2wgdKdXduLsgSK4BrkS5HucGuDZ
TZOctQAHb2l+73yPpqq+rM48fzV7QS0Lr1dvVyb+DkekWBYcUqtcfwarZDkpfqfuQQfg4ouJwYNB
4Oj4VKikzVRCzJ0Kgi69miTt7btvRrGf6fujLwwwOZz0hUZjJMnvi4ZBdVd3T+lJuade+14NRl3Z
H7BBb9kkLhaVQRGtsSy9WNKPnJ21amp33jqUQwEHrWuWfqHpv65oCIvzp70xqfNb1gWezgzazohP
Zd/8EtKoSjvQVA0FcQ3cVbpWYlyoKGdsOX0VdNoh/MeD8P9Sq3AxmHbmfz6G63VMhx6ui1WsOQ99
Br9M2fJiFImdcPHMDymPxCJJ6zPGcLMVF6jIfS42IHAbZce1v6t7DV/rGCbBRG7QzQPYW7XDdyzG
t231LEE3aXRMctRvl8XO7tAON8ignHHRweK/RALxcRHMuHAanQsI1Ov0mKPteBykuH+w57pkQYDp
JT/RjsSruQvovAgR9tl9jEzoKelwreibVfAI6C9k+tOfsC3fg3KLMkxK0Vp7GsKfcL+gtgTKn1Sd
qJoCxXJ2G7X+DcxTrojLQT+sDrNtbJQXIC5m0oZF8BJK7smCxDmvSdq8DAjHyyMf7fRE5TyKprIt
ygBU/3sLumu2q0+RiI4czF9xKh25zH8KLlw82rZCM90ZBWR2iCutMkmMWKoKc1HYI7C10oKHmfP5
YdV41xgtxZB9psUR3trM4wNuYivomYVj4NAIufFs+CPwikLG0g2/BZSc/goLvJlr4jDDF8IHDFLk
4zssjC0251cz3Nn8iZArPDykl7XrADPLgAN1cS9UODNtL3n45CgfsFfobi2yoV4DV1HvwyEwWn7z
Cq+BRGZ+yzK2i/QT/gjwbDHG9rawty3njaSXg7GYawMv7w2nAQNcjRu0iZdYJYyals8cqegOdaRU
EVVaPEuPSewBt/BTnImFLIyzc/ChBqwrlQ7Fx1r7Ezi3nRuSdILbZXDyYWVz1chkxKOAErSwvE3y
RAnjW1tAR4Nfqj6W9y7oEYGuM67srsEe5eSj9cz6eaJL5p66q8YdPi1EKtGPWZI4uwdXikmDx/v/
6W1mk9R82AYFjIGsSoSkVOfW1aBoWlbT5r4krjBN+VeEGMtETByqdz0IdlGrbfmEK508EWVbFwQO
sfJ8ykNrYT97ROIxeilMAuherI9fPY1LrCOVKfBoN2xb645AkfVU/TSVXuYQQE3H6bjPkv0XW3Gm
frFUVjqlcY2MKC6fK+807yu5bitrOHsWPo127W8ZeGOpSOE6jLhZrEUvppfqGh0FZ6JVBgkOxO9n
C5zavpIP+mtUxxcbzM4p+ifWIKINKFNikXQOw9j6x4ofSMsFioKF6oqVFNsMh25mqeRQ2fp+bFJH
zm3eQjSN4nBPfnicLv4zWHcSNJvx+dNfL7UiUu8BPh+y3z+dEo4XEnhcq8phVZYgIMkdILIMXV5Z
VHrE1V9b2eJwicpJ6oYi9pM5YdkqB4s4LxDghqWC7dTq+PXHv7RdLyQ2JRfV78w+/z6nWaTvqn10
x80AYCXaeSB73nF1qeJdLvRHomu9ToWohAMI25cyjjoGmwZNSeZkIURwbBLA9B4ihqn/MtCjovsK
5+ZTj/TK3SbVPv9dnc30r6NS0NM2WVVBBisb6qnI9ZqIHKgD7VtLW59KfSDjBz0C2T9ArD3QCZOI
QhSlrU++80XyAlbTRR0SI18PuZ0Y+IdNi2phUhEgsURIlgENZsufpCgylC/Bd8hROuwvPisnb6zi
WwLub/mK8sQZywHT5RoG72PkAh1hxPjWMaX7AO+lADj7FCbO7wdU761rt0Km8IAxJP79EDur/s/I
Ke765uqVcBTPc7yy42ZA2jW6F23/NiMSL2tLCCernF9SuaBQhhyZgZWSS6ZFHJe38kx+sS3qTTjn
s0Db6gEETGNL8cSooPTXNcxQQJl6iP9PHR8aZ4cCWCFsZPOPJmzvFOtfQMmC81Ww1gzj1fOZ/9dZ
EjsD0wRiN/nE7j6hEmfy8+DLJ3HQIg9ydxqcwxXfva6GWFAi+zI5l6mIHqcrBnhK82OLkTSlk6TV
HjBbkG9/S88fzMnk6YYoC3JZKPdPUss54vRTMHauc0yClGnSqqfDZm3QgQBx14+e9iMX9IRKZK1z
awotP5DFoK6YQJFUaVTV+v+rOGHem0rQGI9QuHNyRb6shWuXJHsHqkKuNa4rsUQDq8ExnjYDwxsW
hYJo1VD4Pw4BTnCtpnrTRKXX/vx6vXhCG6wNOmCiq4P85Ua63g3P3+xAwh1FQePpMJPg8fSCakjd
O+keJQfPL/BOX7F4Ojs+SPMAhJm+yzEFAQcQIZQHflLnbTf8fCB607YpmAw3J545h+NHHAx9RVQQ
7NtaGuNsl8wS91M7p/2J+UGdCqGDWF+RZ/ri0ilEdbj2kcczwiNIb05rzUvI/fjTqrCp1n5FanAy
7t6mBvze2Kqo2Kq8AvjgNvn365USsjqfi5GCCrw4pUvwI7oQRdcnzqSFGacSTQX8kRJYP9v+REbi
Dhi645+wNs8CvQO0qkRVL+34Mb7utFi6hlHAhY8NZwv0Sa3N3jPBk7kyRN+s+hk4vnF8T1fglt/x
CNGWkL+OTSnhgFILWOKMPntEbIeUwiYreWIkyPG9yFv3LFTxG1qrEE2BsNwj29mcwHiOGzFOWRHH
zfT6nQ/dIgel4uDJ/xz72xcAM3PNQ1+Vt6o+E55um18TGdRD0kpMYDtyna1jsWlyTYRd8CAgphj0
2cIlLCDGvjiVtTQrzoRbn2E/A9+WcDjwVDmu6I2cy7DhfUvjNEd7+NhMk69IEsIX0RN7MMNYD0Qv
ktDMk72RuMbzM3+1fcpuMO1Gsq53uVeVjZDUn3qKlCl8tZoHUM83EhsYGgEPE1HbUhUMr6oNjoy+
WnuQjb3tBZYi9Xj2haTIdjVWJxo4UjndnXuPxrtcBXpDZmYP1oLSjwGNAveCSjmgdfV/GK0xS6qm
En0rtIYtQN5M1Hf5zm5C87XqdgQY5FY7sREA6hGfqEnfTEmMndKLUpz7yXUqEV1LXNLMv3Y6OgY6
8GmgrnKEaMuRiRLYcU0/UUU/scxkjG6yFEOvmy461itm33MPKXLPLcI0bC9Lz0TA3KBxbomIsj9f
xROQIqchL1Of1kSMOZ11DDaY1GghsUuB6ynm5RZReTYU173IdQJBZ8gvcoXFD79dW/xSq02d7nSV
S1+OxZLNuIEIw7WBAgPnQvFHJ/JKc4a+Ix49gJ68qkR7uhFnciNUkNHYkhjDAgOgYY16yRjo05PG
6xvjRW05vvSCb+PDa/kFGQkG9eLM3EexnIi+byudpFcWDw7gpczwBODPzzdLROAgn6KudURSuG2f
mFm5eWML/hVaUELMokgeCge5IZ6Y3uwFNAswFkpxevVCpfiIOitX3CyCI2L4CcoE5gsG64mvCoUs
ahcpeH2KaCm8/yw1gGl32JWKnf54kN2pJF9QhoLfXQkjrtyrbi45BJwJQL9eitZdVkDXNpKhgVWr
tsuOkh87lfi/syPQZAbMyciEEcuNTibKXKdLxwqLX+X2EEl7+nDCrWHj9ifNIiPZiCCFAyxcIQhZ
K9H5+IoF6sBUrCoyll5c2GdA35PcUpFp+oCSTB0hyFS4q8sgth1JPkczI8nJdEFkyHkdejHc2Tt5
ykS7C/0TfxlWGllpwIHeg5K7CoaOSokRBZ6nB6CTVtRPKZv3PiIJjw0uDuSpcbusY5JKiRwb/Hq+
5aDs0zxF1WtFRjbKTW0+gEW7CKUbFzubxg4igEJVRyloKKJN/1MiifWt2xJ1fsB7lnN9l+wpOEcQ
Fu14vu7WiJYf+MXBB4Jt2m3bh4QO05+zeCMVpQvi1gUZZNsjHl5h/zZzGWkSy8sx1zp17ZNxRV5v
TvO1+3pKAY6dpeIzOcvvTs34626RH3kReB9jzP6NMKKpam0k5e7hsRIqqEmeKtsDblvj1Y3wNe9m
DEYCWso4iPP8154uFgnaCrKz9Z1LaKhSN5lsc1h+bw1zIinR2hlN2+Of0FI0fOw/9S8l9Ufs7ow+
c2S/c4ADKZaLIaAiKgV1o14z64TfelhPJl0ZSGHW212X7c9kQL9FWN3O+7l0x/IdzG/EDjirHmoT
fPo+QahA1xtGznEyRetaxU1SYGQCi9ykpgmpSjH66GaeJ2AWmJlPhO4eDobQ+ayJtvt78F0mNMYS
dBfDUokXl7UC4Si2dvjmEQ/1SS6RafkclqBJRPBnTPhci0T9hg0aN2zkXr8L0R+y+YBoTmT04J6e
+DkrXVcDEyqChsN0wsecSjUDogfXgC1l9QNv5McTgtY2Xvu7WIGkZjrPF4OSV1W7DSpk713hgXeg
6ueOjnR7xHk9frHXYeDYkf1ldFdp0IjInLLlEPnQqMp4j44z2NAhwFSDIXeSf6NXFj1JNkSoV3ro
WdT5/aNA6xCQVjRt0NTn62aoXowhkkeA7xq4gHmGIK8VdSVlR/waJel/CUzTjjIS8Zdqjhs2R7ID
NhRVv1+dSP+CxAtDPshHa/k/Oe+egN6Mu8TeVLJ9XR3ESQZdqRwB0ICBNkW86jNgrEVdHgzxhe/O
5r4IQCv8AD+3yjQ03mQdDLRZUXsp0Iylkd1ZKAbB7MSQVX0wZnV6nshAKQR3xhvk8H7JtUedqIaX
K/ly9uAf8ODpYHGdFi3qnqunGH/qMeroGuV9FTpGzOeLthH3AI5pZJ/bVyH/ogoCLcaVGxg7Sui5
yyvPBAx6Y6mUZWXfWuXNL4wmzwlfw3kLdKPiSGYEOSRnfd19gIZgMEf2b+v0qfm7wrckebxYD9nk
6WvYHbFTxJQLMiZSJDqZadS4mws4zPc4FVQ5cDLOexAdm7uXPimGkXhtWieVSsPayxoCTHwyfV/o
bOse93aAxA7SqIXtV55i9Sz4/Au+Xes8eilX3+ue5FHglth0LBQGXW7SCpFMyF+liEDssvv+KpnE
+7F+1W41ldpD8uJZiknv6rpSdahnaoOHjo2nhWc+Fc/ZL/521C799sXzidfnhMOnMcOJsYtSxPGU
7o54OMJZun4iJERDKvC6hFv68QdTP0XCW4uFTJDE+B8gVtk1bV7JIsNqWzoaiRpEL9PQ3C/s5uM/
jJt0MeI7oA1s3z/hVpU8dwqT1yKRVJoFBuUo/e55CHfZTQXRMaF6gad/IOCN/hihp1p3c/sNkKkb
yOOXP0C/FKKSGfno0wOaseIOgTAmGGEQtJXdqBL2OyIE/+kBjR6UBw93MIX3SmZhNILfkA4Pje1U
SohKF1b5txhoJ2cmqOBw70vQv+GcZ65ChpZNZ0r36I13F59KUTYZlxIYqNa/mbsgJ4JfGJZKVj4x
jY598BM4A94pG278GX9qrHfhy/uHogdMSxIvLutmg2wdDu7KYxpFWZdKQUN3ipU+/k9AhyH/JxFw
81eA/OefGuzXWHExxth5/4lTuMgBptmsxeuWDNmE+bUp4p17BGFG8ReUh1cBklDPSjzoOHa96aDf
apgh0lvEe3Z0dRst2Ze0rtnhyYBvxMJL5JngGf30mIglynE0G1CZOzQL57vPfXetONTcDfaAwb2S
QDkVGrOSWwLh82Grr2NQM8MOvefAcbQnu0VySlzUuexfrqGGbPb6kBaxLKhVkM5EXQ/j3WlT1g6A
eA+dF/W/y4MfnVTBwROPsPNeKQ4FKyNf2t59wz+5E0WMR/rsKJ2hZYzZ//wtsolpKJt9glwibI6Y
vst9PHW1FswKQmXzWLAU58Re+DQuMgc1U8D0NCCWmKwBHPmx+KilSTFTq1ApMVtoUxdBt37BEFRM
kzRLzIiX6vAfgdFFeqAzxN05vqK103yDvbTTOHjQBLAuQa6i0XciPkVt1xhZRLw+v7dk03Mjg8xp
IGKC8n9HrepmA2JGwSyZqnfMlcraMlfDTkosFfe2+bTKJb2kD5irETWASUH4DzRmQK5rxRWINleh
svCKF9xuBbYBxe8Py5Yz6/4nEM4DVxB6l6vGZR7xLhsUQhxV/tJBsA9YWg9XLzxatAoB5ll7TUK2
zBlPzW+z8c4dzVRIeKqmUBfkR6buPv0u4n7dayaBIkD1zdYW/A56FBANURYlFZZhHAuUV/VYz0pE
7LmKNSl7gVu6KIEpkrWf+Lpwl6Pbtvhkjw9V5NUR2wrxSnQx97O3LoLsOG4eL0lGJhPlv16mb0/q
I2ztHMugRhpZ56zsndiq0nE9YZygrVZZeazOBpFH0yVkFyk7zAEUqHR9pVm3Wyb6uGHlpWwqCDCA
tVoE7UOdfkmCtfxXFy22tPFod/yS6cRw+UD4gpxxVzkAzQspb7uTU54RxIOSEPn/bUzvLWjtivxu
rePOGzMAtj9kVsOeS04wbgBxImpd0NVAkCDCija24RqWzoQq2kNaXSuttPTuoKN91M/p6gUPGLrd
lIVXg3DX/4VFivf8kHs72XGQf5bqHyGFEzC4RJOrJLU4mQ8vaVQWY10DdEMsBFgOaWaMwN0ebyiJ
wddXxzoQuem9jDzL87MCPhar+7OtDz/icb+TmALwqmPlZswIWiTwXrNn18KupIjgMyPUySxaTqed
QewyYXdanhR/W9mWmB7/dWRiRSypg4bi5bFKS86Xna6kyrbGWSsYx2gsQ9oDocI4BIReOEsXvKDs
afSx88ZDddB9UbmLBnipeYMfQFdelllsSGcCpCw3K2NTWVD7HQA1eziWTnjn84wgiJaw2roG/w+b
fnEcvUrmCxQ/4bdX+nTnmV3NQLwaglraczDVJTo6Ohsl0LYIeFwZfypv8sD3s1/3UQ6lkGDTjiXA
qyQhL6BjLxupd0Tcx4FH2X3qEDiEUNDFxFsc/c85aYEzuW+m2youbgV8K0Oum9MTjs+vozN4PW5o
Euo1Q31OE7kTB3XRPamj1jLpWWs1y+u1p7GOOmjcR9U98TWmqkRbPkJmwZUVhtq3SVZAqHyK94ea
LsqsWScDvYH+rYJsJPvHcUrF51m076i/cVd+feFcxookhA/1XLYDlfEUjmC4b0PQkdefGePmuoi5
evu6di3vtVJ4MKq02LZVu+PYbQg6FeSlwi6Vu3D+6lSb/eNtAHDD+Msu+LBHV4+DA1dI6sWXQcLY
yP9djh424P6MgZCmIJEde1LtOr1EeLOd2gWyrxpjs1LMCkpX7+tXpQ8lOcCoHk5cqI4B+pE/yJ1p
0SQZGYH8HtWBkQi7gNxfgkT0AT0Sla1B+L3l0zr1RBFMvAou3F0fOpgWfexc1dAFtyVmZzbnJrvK
rEOLCnW75FNPTdKFAGZF+XRH70lKwtdFGx4XJcQtx4RFA738JxXkAZuOF9ycZ/vEjIKJN6WtHEbE
pwps7HVVfXrUuI0YoZqcnn2dUlPbacrqgdOBeKQF8FxjXGKZssAekD7H1hPQVeMMnwLdAGcP6Nyv
8K61b9Bi7BdcXTIqJoDBgFQHMEPs6BPd/ZRZAG4JhEjCd20oPtF+K4aLOUcaG9DP7O2Pa+sho4nG
MMwS+kLl9oX1PTy2i1vKJ5u/OkFG9eW32OfcyG25NAWpYmP6ZvteZ07jrJevbPsXV3ykfOLnPxCh
Vqh0LINsGC6M01u7eXdPmuV4ZBDGv+AigclIlz1zSgnJyZvnauw1o1uEIySQ4KEtAyN9xx1GRhZJ
nOcEi4wFzdHj0mmm0lt15bHOQjm6cG78SnTjjgfhqUAVH4vQ8Ww9ldKlkM6q+tfyVPkV9p9eS3Vh
vqIlBt9NaTWaQH+dBZtVslYVlhvzMVmqjxnv3LkrFX9MAMPf9+PGAZ8IRsqWc+nGhsmPBgIRaAzV
9qdkZQnXJUhbecuk+7ksnIOxjuXK/1xhB5jhiVAsJOufT6NUr34iPu0xc9ue8Zon+HNsJgWhrjNA
SkFb8YNs3Z4RATpERX1I3hBlyQGRKTivwSf+pYyFnHEY8+T1BZRO8f4uanOFFQbWS8ogA7MoFJqu
Eae6Ug6VWKgTfO0Mlc1wcHpbdeabu8O6ob3Y1UVdfrGnU4/C6d5IahnOkVsFUqNYFO9VJvMswatj
HYZ6LR3VENa9SyP/xcHkfTyq03QBV6mzUC1pxitd3OBzvsKFOnhEzEuPWiDVyjM/jIK+3/B6RPck
dUEZq5n0TkADs5zM8aQrU8x+CG1vtF9FovnYNyAMNkZsU3OnnQMkvNXGD/Xehikx08V9n+/VMkbK
kmrUV+2k2Mp8ZIz4k9FI0TtZp6Z7S+O9aCUd26ZsO+/Sg2mt4PAyNBPGpCvfbSHigcZb5flKA+Sn
E6w7CpOtI79YZYrxgLHdIv+r+QEBWJbWxt+C7HuPD3ZZTIvH3WKBQo75EdBYMBaGFfebPRZRYI+O
CKXa6fIZMrToqADhvQA+Dsa3c4J3kvNJwQwvbKy6858PCNV6eDS47Kni88pDak8iy1zXRI/q1aVM
yfxGAtRQXErLiRFS2/Mgs3T+7q0YlV+J9flArwbSFtUqHUNTLDpRJ72xQ0/1UL6eqpY+PvwyWz9a
93N9YzX2wn27Dted+t5I51Db2/fH4ZuS28ICnUp5j0n3u6a4XHPmZGiZZJctX7Jrl2VMxH3g8WPe
Fd/WnooFevPWtta8dJOKb4u68cbHND908LlSOpNnkoC9B3e2W8PbjJT2my4LVVq2O51UH4mus3Zb
fzNzzhAkIbz6p6t3Ez4z1/YMKBT8clstZUBMeA/6A4DHtEJ+HuC3tVJyntumkidKKo79GulZlIBs
H68ur8oLgQJbMh3oqN/dXsuXUbmqvXvWXVKojsiU1PS6Ezq9MRwsogKwBJ2PlJ+NrM3jUSnhhCTr
3tmbD1WeUqsDoX9k5GQkeYK9ASA8bxfmyu6YNlrMnTrWsmZfZjo5jx+kmLKXwK8OpIGH3sPtB3wp
r08x8Kq1NCPdq8wl0hGXrVazClza3/HnNQrByQfLJm+EW2rphFuXxYsetMZNZid9+rw3uqQPdm5F
pU8J29ZwCl5m3oupfbUi3geldrPDOUjTmh71RbngAXjefDjUGeb60vTzLo0KTWyrAVKeIk11/2oe
wDXznCB82OEDBZGr8T8SNOM9mYB6qySJKGGfw1lsYv/WA2fqS4a1kAECa/P4ECB7AlSR1v1bZq+S
fSiPAWEMz8t8XNJrtor3jYJaU9f9clbcgy6fLzawHGCQKFkwsXOsevT07uau+Re8BwlIIbYj+KQ2
5k6vagGWYJCrtCWsft6jDQyvDb6q9+2xqff6SzreUQ2LqohBmPFn1Okh/heC/RyTJylZnrfcvi5N
u9HA7S+Gsa02Vz8pgYmJSNLA8Rdey3TFDOyoz1qscDzjo8Ddr5tF0vkYksTiOHnizhB+AZn2lkE4
OxgP9WIoJi5L04eE628BI1v1p/pk4zl7y009QwmoqBnb5oQO3nWf5JPuoQ/TCBurguKe7bmvPDbw
mEb7a5vtdqp2JSeeTV1EDpDkBGCP/GYcSlGIVb1qxE5BLaFGJWZfl5LuXgRLBQ+ie4e/vDAh1nUM
Gi5MVgt1lmAt91TiXdHVwEWUOlGY8SWNZD59jkcEqTympWYprToUaE6rioyWsFc0GRS+fgutbfJv
Ye/kFCyql3pj6iEBjGX6icmcaJyL8wiBvzYAw7kxIhuTKxsb29LccgvJ1oBRCrnSJwNSr/fimcBD
o5lOjqxmNfDeDEXdGy4WwdFQBk+5Arx0FfexPP9q14ih2K9k+JE3Sn9GLzLFQiN0pooe2+hekk/s
+B8tJRHPOG+gf8og5kIx60p9NTzD04pGNjEAq3hcFsn5kph+GW74GXPp1IOfj/WHwQZ/8ZsYkPrP
8KXQmfmrRQgFcJ4TOk7J2rhjdum24bz3xKeQWHGw3mhfD0FMre2ugIZ+XHXRltoTz2OnRDgfx/5Q
ZB6xZF3vFvMhckztolUlYNuIkbnvT1aXVtgPvYVyar72JoeIwHZ+kOuJFpnk+tOTDKz4CPXDWTbU
MxLuEBHYjaGjP4SZqbhh3b6XUQi79WiBcg/Z/V7azIXeUbSpQVv7zqABfkCb0w4XxskU1Zv9+BCB
hqZbndGG1EYrMuu+CRSXz/sH2y4jzPPflAk1LfR+VyrisVGfIgZC0QGjVK8L2r2jSzUbyU7oONQG
3ou6K7fF/0P2/hBORSGsICVapn+aQ18tlEu0r+S6mqrix1vB7Eg8h8OzkQVF90EXpLrRzTf55f3g
GPdKWPUWl2kmDlUzPPuH52r+1MnYSjpjf5CSaI8bBPlStIdMrvdI2d+0R7CnwXLk5+wK2mQMJIn/
GMrBC4W5RXsX5DFbwsw5KICpW2CUSXObHkIn0OvoOatWVyTU4DfSPdxJvpHIZQ0mpF4wSCZRGXBY
3XFMpnpuWn+zfhAtRea7CDqJwByCNA4WjusX50/brX7jVHKG8Yh6FBUV1lt1bWyHSDunrUb7aJlt
k1ISY5Q4z9/Wk3NHH2mKz1MVgAptdUT9yyLKTZ7IVCrPSCIIc+pz9m1Qi0ivd48X5Rmbj1s/HkKz
AunN1MwSOidS8O9dZ6SgcN0ONsVaUGXNDt/WkPoPO8vsgc8mBvHGU+TPlcnfTTyGvwACY71kAIZu
Q5QhntAoTtAk6HJJU3SuzA9blqZu+vRzdE60phLHAYv5LTiaKTIv4lEYVPJ4J7LG7NS/Rh/LAmNn
TeZ4u9ln87KWQMd2fzN0oPk+CuZnGIFieD9k5YUmjthrHGjrDmm8EYE5nDhv1MaV7vp5O632iMcL
AasvSzcjKDZyVrAV5Lg3vRpkiiV8wbO105bVHOKL1r6M6hT15kFlocgqiWH7nIhzytRW6Jtunf2e
4vnhVtc9m1/PhqaiZS9WPzeCazreSDS11A9Nkqyw9K3xycviX3y0hMpCIK6m+/imRlofQ2M+JL4u
mbIEt7JuT2vV3viDVU9/Aq4XsnuNvOtDMO6JMd/JR672URE2tmhz+fNVL9elJdpjjgmKExabuxed
ikLXnZjgFIPOMT8OLA/cidKSTo+6EiSNtBRh0bvN5VEcoHjqdAgMUJI1iwFdDz2Y+MJyqyf31TiD
8fawQrUm/QVMa+JRoupYAonBcJHpFqHNf5fe8bbTjSM1YkFARwWjT1JIviXFuDMAykhrRbkt6Mx3
It2o2QejqvqOr6G/4sA82cBc9CNyqnNm3nDBsEqGsm/pVKjXTzwVhOQuPgKxmR4d5ity9azAkiDs
mcZliFNqh1sVKEXSf753pDvtBCYEmBxgg3lv+SmZnm/GNLC/h3fyuVhD6KsCodEKvq2pmxnAnoBL
jI+EwPR7FQf3NHIeTPmDElVpyD/3B5bSvePBfCEXNnl3LCn3vIPnvxm7wDBwW8bNo6dAqmI4q7va
YXev0Jg4yMtxa9Rb+thjz58odRG/asMbJykSu/Yk1SKsTvt+SsyiAK+LGhSUMFI44lTZqtPVZ9g7
O1EgVb73PQFs69FGbZZN7qHig6DcbXMQ9541jQoX0SyPXSUiWwt+Lz7Kc6JiYLG0rgj/4QetT+oJ
+/R/VmvqDyBOWgkfoxT/oJAIoJof2iTOenPSMbKzAPrkwJbUgnsTaAQ9zHRaHNH9+QGI5B+eMrxk
f2Y+eP3mO08kMfsntxLUJ/17WvC5c4XBD160y4Hk/j3Q6RzItISBcU6r3dj0U7B+twolMAMuJ8qf
GC91JocJQeLggg+k6J06FYO8mZwAoUf5oG15ZGEYnnkMp4zvHnGtiegveJBtquH6fyxwuOuMb13V
g9MvBgOvRh2fbK1hhcDldkdRN4ScoXg3qHkvwILXzcpMRB83S7qbPGdvDqQl2ZAGRoPckWYwPEyS
fQAIQ4Ly+OemBwxMK4Xj0x+XcCrF8zr9je5LAh/OOnbH+PD/S9BF6fKfIGHLcFsqYoquWbJvS2Ya
4SVL6fZomGgyWtPFl09/goU3nkvTH4jMZur0yQBGTo+C7K0klDaTuCsH/GsVJ/oOkM8ACFthOfF7
X8I4lAwh1U7amgRIvjRkvlfTqn8EQ2HUBhivddLhM+Vwr6JcGPUM5t2esIltRJ5EFqpMuIzJ1bpJ
ddW4+fQsBJ2WFPV/xxF3JKK0BXVPbQ5aX4j3/WQiFizN3o6dw1Squt9+QntiL41FJBpepXuNMjHu
ccJEoDRP6sclFZu7P0n0gZ4IPMHGNu/byl7e48xSV5GwqimMtG0EHDq/NulM0do52NIS3/VZKRue
c/C59YpR1FINIaIu8uXbmKWfNIrI5HgiweYC6muoQ/kTggag006TdBQAyQqs9euYQRrXKDj7OEN9
5JYi8rd4blxRpkL1KwFnNkOeLiwFWN+YXjzC8irHGURheDRXaGwULzCnAH4BagyUIa+yzJ8H68So
96+/j/f8nEXyvW2NY7pSUu9k2srrw9ZkTQfLwNMcObeWuXhwoVyZhj2EndWBh+nSz/rWh9kj2TY0
VebHBHGjgvVmmf2lqEqB/Hk3p8kusg1pD9xFXD5a8cmX7/4qISdsPCORxcZm0mG317RDeDnixA2A
L9VRw8CDOsHhczUsCewyg8j/9/ALZMon39A1rbkHPx1m/Shd5Q1fZJ+oL1zFCz/Fj7qvpOwZFk79
mSMI25ceyaAOVKN9uy914wXRrBDtGnFQfQbZKMmBN4BlhA8zv5yarpdOl44jItdtpv6NymSRt6gB
0yio/1FrWzjAhbqNiOoMtKRbshWRYLgXoDREn44nnUAoEQigVGt9mfgCJYpK68Bh63f4CZQ2LyVw
/dH0IN2BMj/2001bPT2+MLGDcOOahBEZmFspO9kd895TWfzhLkYEsszYgBu7iCmxmR9W9cy6LG4a
sl63LfAB+KROBvXynUSymocA2QGEsiw2B4ouDIOq3GxCk3s18suYcia/WGt/TAWzcMh02XIRGtzX
gGPm61Cf1Vm07PZLyxV2EZziU3RU3jShf18kYkR51PiG+9+ChiNi0i/B9hv4A0nlRvCiYFtt/u4y
aJLUl6aqz+5p2Eh7DGodpT2SqcoP0l/1Awunxtr0om1qdevC5BachZzBW6LhA4XjcVkjM8BWy+9I
Iz0UD/BCpSpVxpQ/jcmAEtSLSauSUoKyG/sVsVbLQFHiaEEpBjpm+r+2pkI7D/YJWd25U1gp4BmC
4B0PQIUn4vvYfOXInDO0agUoc2q/jFPca+edHB6SXxnXtHDwv2jOY21CUKuCRU+9l+RB5e4FMiRD
WtqQnT2Lz4nOhqOLjdW4WyGTNG6/Ku/oXriq6jbXuhWArR+0S5XMeeyudzNoLchdYaPruzm6EKEI
92v+obI2mxub5df1cbLrZ5WdHKAXelyH37lGyqtoLLj/gWQeE0fTDts2ml6tLnbUg0WYtXMM8oX/
ZeCCly3aumBOgavT3YzlGIBa8oEnBM9dxSgUw38ugpBN+AFfqbjuPy+95QmsPdy4/r4vtGuRY+26
Xi4vZsNE73vjNQ3cQIYT5AsEGNDegZojs9XjQ3TRFoWHOoXKEHdbUzdZj7nt+FGkj8vq9R+oIKis
T4vw6XsSUB0mTWAme+MIxwmW4tmwRQM7Gz3TX6/u7/6DY06ArlpVMHnzeUkr+iKIqSHxsgRe+EHc
hhWJN1Y2oHylVs5KaksOVobQ3L4b7BANuFhtjPD3dyqDla4l/UbpaJaJPOYlEpb5gY38+GbFymqb
iJdNRYfLYv+/25eyPDWlQ2tL/NqyRr8p3Zp6lu+ox9RZebzr/qX02nUQomIzMtyVOBktsW6jzxFN
nPMXJb75BfaBNzc50xZ/OqgyBHib0y/sM0OEKZx4yoV8dd5tTmSJ6zcD5uFpE2TPFK5aJrxH91bk
ZFrV2JgsfRqym14BlHC+uGV6/78isMl1kQIBY3UapLse4Wd4aFTxVFWpBnAQ+dO1PlvBLf80n3bF
M63AhkwJ14z6+SLc7VBUFv7gftK41uqY47NqYDedK51NBp+dc1doKx10YCW17sMaH0PKXmBYzDEH
VNIETLl63VbLSpVYeoxGQLzEtf7nVUy07q++unGSCXKGvx1wF4oMhqHOHwWpLil0BhcfwErCyHZm
uQgBuongvFWMjCThphdC8NTnI01N9S8JtgmaKuvvTB3GkkK5139wh9dYGALKF18nYnPbEq/DWQ06
8CIoy/V4tlFMv3mMIcEBWke+a4wpv9Edjof4iU8znw6gFMx3JHi7Y3m25W+bV1KuXE2BmBIkXLdi
9h71LCUNF5G6P5HWB4+HJQuMbsLZ5jDpacQmu22wSl68H8z4vuvD9vDqNo+aUdqNfsC3vOZYi8ww
04nHT3O5htjGskA6cfFfA7JFXdHyUDxLQ/haqZrW0GNh/f/2CegWmUSjQu7WLSNho0YGXAyNVlCF
lycmL4Tyf0upJzN3IppmmWxaP6pj9tSjDpHE7FqVZvPHLaB5iweUXhxrNbMzm+35ShBsH+XGJXZ9
qnWGAHbZ8PxsJRsl6EnDN/4PdDOZH0Duli7UZILZhOQr8JAC72YtXXoU8otK99DkXBL9DkUpTVsw
lq+721QBuKCrXwLSwTBrygCo/Hajho1S/ZqlDYcKsNVv41+63NFWIYVMRY9M2kF1wbhBdBpb/D0p
3+kall6iDGkCNyyJSjETfxHE2UEhA0qewcFXSBA2DNSJvzbhc2jw7X7qk64KrSQpgvqe39w23xwR
9mtsmiuHuDgedpAWReWWUKMptDfMFhVtKTlptc3jay6NCGm7yxjAQVx8n+DAuKcrVrHz6zZScEmU
Hgl6el3lmVsNkGdmEUzVUumX9bH31BkbJ1FsFfKxq83BGKOC8jsUP6Eiz8Vur5amlob6lMA7peWh
aO5vk9yjhuMYzGVN42L48Yzgh+cwGNbhaym/QVAxTFT8No0JQaAfYkTQl7y2VBAPe17aqZdIUTlR
+S7roMSLPw7ji3+U+/th4RSw6W3jkrNQSl5G+jdbx25JsH6kkkFNrbDNbuFRFiHOQCMrwOslwIsU
uh9rfIu/ShF/dYyjSmWGY1u58PqpyiCq4kThH8z1utHsx1MSCORh2lm4YWpFJTVxdDQpU7eqJP2i
/HYf5yFn546wKUgPTeL5+BxbTWUdnhEuB2sfZchhmP8K2d4oW+ICuLt4gRYHDH30aW2KnMjOiUNe
03n+qm2To4cuNDnxiYINn1O7JaAX8LPuQPYCvIggK7THhjz2ESkN5zRXzyZ3q9PHBOHGrvf5/pqt
BePgy5KDsmSt70tIx5piIbExcXAWILb29KJJbjNSm68OwSO6INUp9ykvryMX9MPno4xlkKD202ES
JuCXbfgu9mIFMWWPD046BlgOl3PsonbJDTvPPa1CyYtE8Hx+t+4wPDgDFhN71T3XN6jrBjs/+/oi
IFk+p9j7ejNgH7QvPfXYVMq5iCgo8R2jrOMIscMsRETPB5wb7LVqdqxdZrYcyKPW607ohqI4Kmx8
vJbzHLN9xXeU5saWjhwRlMwC9NWwm8GEo5YoAvzoJyc3pFCkcxnN9T0/118uCCVS6tOWnRZ8bppc
5AZglsHSf8r9FrgxXfHPVSJb9J96AfD3D4x1paTduBW6wq8VTehbFLGE7mvIoQu5G8zZjWRpoaUk
x/B6I08Kix9mxRNZHuNev6leHl2i9F5CMNWL2nRlUeS+qGklCu6JZFDppHMaeyr3TjDPiP0Xo1Za
2Dqfw1BCh2kAdlnQMoDsC16+7sZyK7C6PJrLYBzB2fjvTbLZsW5GLoEy7fGgCVMOmhjs1+5FpGhl
raE8Ecu7VVoI3iHQ5zqty9FPzL3jyVfR051xUrsmsMAKMSfhFFCI8ZNKNrHKn83HSPbQRcAcWmjl
79mPf9EUDiEcyHHxTbyX7tLqrydh8PzB+N/gmrwlgOnPScH2gBVElBtM1FdI4x/kcnZsKIn4A90m
GB7DMdzUApQesR1P8bEZUJnNiR9CVJdx/V0zGmQ/zjqVmbkw1WVXmWHAz803IXHy25/JrA8vO/jT
5/+V7Dh2xIoCCBWjJI6y9vUhvIdVpRQRtl+mRUB2FzMuwHtIbKpjki/wDjwOozWgRvZufGdktz97
UWHNzkU4Yx+NsFijmRZA28GNwhXqahU0fgkHJFxgPM5TtcOzAvF3HO0jCl8ZmIb8BYmd8oeRiKPv
W1ZvmTigvot6aNPlvNMf/JIbet8nkNodtkm2ilhiFxMpi0ilgwI2xYZCE3dpeiw389F1fi4K9r5s
PteNz6oyyIjcGTaeHBTvu16mR4jJ4plkKRQxCQ/aKqcrX+nr26K4qOdukc6mRNvhnckKp9643VUK
cerJtlFISjUJuz2WWX9mndk7IEvc59PFqRUzAOaUvtz3QEATS0hpAg5P3O4tyj8f3mvqQJS1OVcV
ub0zXr1mpPO4jJ4V3c6YOLJe4vmK4HPqJ1+UqrzKCOYiNPT6JLxHz/5pGuRgd6Y6IKO7Fx2BKOsj
WQXZxFTgNEZ+4ELr1IxYBmoHghUK3qObGDxQQxZfakhJwbV90D0rqv4hZEke+sJg7SxUMw3zKpYN
HZVkDRSr8xGDJU6PS77H83rnFzCTmFwbDS+cLiaKtRuvd76GoAeaV8kTw0yPCKu9ku1c3lGkwqjN
xtJqp+qZag1/MNQgmZ5Tcu7HIiCycxezzdNfRS5xCJE2BLpw0G2sJUREIkYDVQKV6T+FXgz/mwEh
yplMLH15wqyzZZbLLxJ0n4FYMxhC7rT+uHHrhXhz8/IkuEPTyY8Bn3XyFQJlTRqc37KvRj9zqFBa
9E35IJ8Ng/pICKvufQ8WTy6z0JZHeQGJxS1ZIz3YNFWQI3z4j2Vr1oy+qMsN9+MevTB8KrSpyz2h
PVhJa9qzsZ9oSJ2/lOsA3vCV5d18OqQtyRnV3oTqHfUmJYUyOYZUuaBVSIrSQAGfo4dEOo3rIu7q
IgxsxaGfS0BxDg4pEwL/s8j8Qc5J7drhdmcj+3/Gb9puVYnv7KqCPGqe9zrnjkaHIx1G5+kM+qk9
6YUeLHoW4bg6iYX5MRaFTKKj8wEvtLO888f+Qdwxy/RNnEZVhFDnG1a2i+LiVzLwAWRX03qMou/I
oa93cZhMO/5uWN75YC4sawfnx0XY1yfbGd7gOyxk/PpcuSMZJtuEld1fou9+kzTgyt67N5qRBt9D
1GUHCUyoIhr9Bd+SrYNVb29xJPixFmNyeJCXI2u/FXMWzVf7nS+epNoztMSgyQw2kpMZpKTUnPPd
bg20sejB6nS16pVO2UxrPZCYR0OuTFjL2W3pEadSttkVjmodIb8i8IKJpjDZfJ99Oe3t1s7I+992
Pp1AeAgzXoFve+N1ivmPkHPTKlv6lmM+EZsE/Wfcuo4evM+UOhwkCOe9Xes/jtvkmHTMcvdi8Jr/
woZmasmUk00hQRLYJ4YZKB+ghWCGy8rARsaw1UhI29bmDGgFlRGCC20/7ptk2SNSkaLHkxlH9cbv
rO86kildqjAGGBbBh1B1ycPyURluQ0joE51mF046c/VPgjhdFKhq2sAE47uC3VDS60wkIhranVEi
FGoFK7s48jV1bXGNy57Yewbq6k4dGsL5ZLTVw7uRxvph3kDLOUYzPrEZiAskrXtXnI2+ECgTl8dO
2hAhLcIqTP+E3IVDZhyMPWcCbku1esFSbeaqEOkd3SBXrVJ30h6d1kki/8OpjypZHkKJtgEFs8yi
n/J5P4qcJ8TZSP9BczrBQYyFu8FVUMQV/5U3dcpZGH51BQCxTEZc3G/0o/HJpXHsN1y01a+XBW7s
lIYhJrMxItDW8OxoLalaFglQrbpvXhJkgwl+s5Nherux3y8h3r3daEF0KIKahY5R+dvh/FEUyjdy
aFJR7rUiSTci9qkWtwGGA0Lpk9HjC0f/WLPVzouj4YMZ2uHDlMX/3LQ4rmr0UVx+iKpBsNxbOrmA
yBqG9zITolJfct3JHIlcUqiyhDPl6gb8XtcyEzuIg94eFHfYRbYco7IFpN3VlQxGbEbiMzzMOb6G
LKzYluMV7S6pEr5i1VeFL6hW0e7J90svgZoSZp6v83z5uHSoSy/zM6PD/VqJ2m+7wWDsKY6qbdaI
7L//EJ2OBpFayHMslw5b5ESO+ng15LobHHj/L7vg/Dv5fpHRq5QfwCNimdXIEuNYzprlCTmNSD3v
SaUb1L5/4MVFAEnfYWvYABIrfGwNGcQj8MNlnA/2Z5O1Lzxm+VLJ9IUx5KHyyweOFkeic2JCvBGs
Se2ipLsrGR7x/hE6fAWHSbHzFSQIZ+NGiqEocu/saYhS0NNYMKAEqhh9EZyFGF2ME2YnpTSNphEB
QWPHowc2dRjOeY3e51dMdurRZv1VkCvlRTAEJ2osHo34IlnlvvJ9W1O8CKq5ttjW/Ia0i/cA80Jw
ydoyhjFEJ21K40yFc+I46dAnLF2gQuH20T++pMLipAI15v1J44ZAon+UT/02dRN6ZIjk+RZ9yMuC
RcOwuokgAs6Q/FzidrctNlMoEV3KtgivAZjdxY+mbxw0khvzHC00vAmsQupYJSd/gL1WyTiEubOO
4Xv/GO4wO5hPiK8Mzp7kQ1mAEx2MifOY0WOaHChFVemlnZ2GzoQkSDit4W8V9nKTeTDHAh313ssc
xMn5h2ywBOsyLYkl9dSD7LmAOhEZlthn2p9gXrx8aQij6aZyo20TFoaGrUUkc81z5mJwgzQYNYBp
SS5+aQUMjQNkUBABfbQG6iGPRrP1Lwtbxq5/UtA8QLOozOu3oJgBm1BLK2zez+6vh7NSrXmlGzDd
ej8/lr4+aW8dS3K7xGAm8y2+6paCvQIwW5SZr/hq84fxcG733vm/H8F/xhkP93l0GPMoNJ9uDx4A
evM4vakztm2V+nc4wTeuGisEfkCXzxOKGtZGUKwMn8QTJaO2FH6qldMgpr9G7GXK3ui6Sc1xHqvc
0Rx670ggUy7W3/p59LLpDdOAMyDE51n6L8y958LEgkKEhuoAYHB/wJEjejTtcLP3mSComH3NxxVJ
LiROHh7LTkOq8e+6U6IBNu4nhON/Nf/p6F0vtojJ2PphmgR90rFX/kKXEkkBErs2g2teQPZEnw1B
a6n1yhBSAjBzkllhZmzVuW9yB4i1+YIIQdXtFS8NVCzTIItTzcSfuUyXg+FyFClhEZ2asnMMnqpZ
ByIIdf0iNi/FXpM00DZd3lo6IyKded3836+6qq0n4VNCB0fbVU/fi4ZMm9ntxDKiBhSzDzgzFrVl
2YKZ9YbCBE5R6O/jkcQ2LGlpEYdj3kXcYfXSkQltGXrWUm2YZC49jdJ8LrI86TKm1IKx9Le6o5UX
ZrOqbbcBX+aSQW/tZ/OEiiXJvuqs43s8riG42lKPXOm0LEXtgDgtP4oXO3nS+t+H3quJqxacQsNY
AEouOPjytkFsrlfRaFwtv0IsMoEQaDTo76FeoNRAdT+Lk4piQVPZ2cf4BVdmWAjJ2JEb9/2LY1db
KV+kC5THq34CsAOvtMS1VbSYEsWxHQ9mnxDhx2oyhPjoQSajbcoQnENKjUJFq6ifi79mlPaKPrEa
ISwydyoEg81NWhGn2vWzUZF4a67Dw+75+fn5CiEhAJKZSnzKhYYorTkTXNxSe8M7MddK4FpTR5ds
1+VfXIORsfoFskgX+YAqV6tDi72f91YzgYxTG5CEmit4qHLs+jgfzRxKfvAF3HXof0X18bY6+n4n
ABQ/I5bFzghf4UdQE5Vl1mzrlHG5FVV1nrH0Q7pu0QsuU2CyH/Af+czKRhPM4kKTwI8pzIzOUink
vLb2rjNsigxPEyliTz5kHNb6J1bu48fxaAecxtyyCu90XpiabwNay2VdRhAlPZ7N6Lb/nCwT9+Bs
34GGiLrcCZ4hlnDS1cjSS06sBpNcY9SwG9Hc1GQ2eiagOziTKNWNSeHKhpQ+EiORooopD0PjjM0D
+oPph8s1VsqLSRh8T9QkD0aJNZj34+t3vpQuA1UREoDP9VGvJKgOyW47fH+GKLiUJkz8bPVmaF0/
T/OJOe1ihq0HUA3ANgh0s5wNwNS/Z87YmbUXyFPTzPp6y3C3znp23E+p+9ZsMXq/wfHZGlo5/y7P
gLw+SIk2Sn786j4W1JlaPoU/LuYLerjvnIwFQtoh5VQ3v/7hJNnWJY0EB7l3KIXa4YEw0cuLbLa5
S9fR3HVBYZm1HS+3h1u0EbYbV70XLw947T0u41SLtsi3jk6yT1fHDtpg02ZwzGA/1pAAYBp/BMgS
+dRK5wBYFU0iBbdAaes+QyLK+pHR6cn0izlwod5Q5ECUPr3px1nRo0J8gG+ypHfOUx9zfdxCS1IX
hiCM3UeNzbSGQ6LOvaZTLxG/OAxdNYmFSXaO1v7Dk1PA8kP+Ya6TpqHq4HXq+f2Hzu6OtgOYJfn9
/Iu+rPxBRJ4E40tk1GZyN6sYohVOb8UvAMCxc/xiJ2k6759jIQB8JxO5ESkMsVIcl2yCA589XAnV
ri7cMPNcAfufM7wydmdFuh+ouWY6YxlyPlUi70Z1z/xKutysfw8vOCAVzgHUIIpbLbZ71V1ADXqj
bQKR7JQcEqxWvXIwV/M4AUlzkdKgm1/FuAL+/s2T5s/TYC+HlnwOOViUClaF/ThkeA/9sZaI8bMi
1uO3rTiCrodEvVZXdcTpyYX8PuJJhNyZ6qba/df6/rOT8EXMutfFoDGJuZMwoHt7nbJnP8gNJ58G
gFIKCnWJGgp9kzmPf3ipeL0cuN5TG8jf7J1eWZqkg0oeAjiVgaypB2vs00ZxoJJD2HuRF+8D6xnz
pNrPYuaW9HEVagDkdMu6O/pLfhui9Tj/aBpfT6BUKPUpuB/iVcgfk8qykEzRwLa/sAPk6KpXzbjc
ix38+Hgrltp2nCCndaLbUMvUw4e0X0ESQpV5nNJA+wGuN/C33pEsq4QBNTNSbX5AXE+w1hhMilsY
HyuFWwnzLAhGHiVGO/AHCVm1ydo8wp5QDzP2va9bhJmoA7DFMIfcffc81vWdc4u1DXJDD9qjGdJP
S9ZMEpONHADL4B8sW4ZE21tJzNy72/KfhfA1WhGQELK4IQ1WqBv9MIS9kTO2yYzzw10bSbKvJrcY
tVBm3r2bxkCY259J/+XdIqzCOkb9DUbsHzei/s4HAAeVJIbexNwj6w5qgNrLTwj7UtlB3J3lyJIY
lygqWLujNDgTZCQZbhy5erWmy9mZhTGSqvoYnLq6NaD0GEqFz5yU5P1ypDXTrDdAtWsZC9CVElW9
5k4Y2GRxMJYStXh/hNxr4LuBJSvtEAgWHu6nFAbLCMiZfYanvm+d76IwZ2nM5wwfZUpnI2jsSA15
zGRtyjdUXopdehPexxOIAx237WhQPGv5AcxpQre1ew/wkFKKQ8Nsq1MEXz8yCEjOO/YOQy61V+Ck
iegACc5ZijMG244K8IIvFNaCZsUOZ1n0l1e6dwA4+2mTNJSjGXQCQUpZu238Qb/hZxenhNZ0t17o
JiI9p3gXDSLFBXuk1bw9/L1OdSSpV2/c52qIzDCNlu6VPPmVguhkgBt/iMO1+1HfwvIdNMzK7M87
iKWSx0oBAUAFhvYT64l21lNwZwVP/kZjv74s4aCaAL5zymEw3a3oPDbltw2Ew1VFeRTq+3jSRM6v
/Q2e69n9BzPr1Cnrr4GWroz/6kwe0ZbXO99m+rvsYorYRWih2+6t8MgpADxcgbtDaU5DD3MogeXg
OYxWG9ZLOaFrZrTxw/+eFgrCSCGcZWcuPC/gaUNow5biY/1T1tED6QeQ7off7mkiV/+Co6ZfbG8K
kqCicaP+Ga9gw8mtSRgHmsaEwCYcFJ89uIeZJldW4WWQPVNL/3elELECbHXpQQDG1aCfD/iKqvLw
C68DXR06DnzBMzf+TIwSHCungt9YsE1/88ZBk+wbuxponmFeeoMv3GMvZXFlkhpwToDw38XW/HsW
RIcWEeLdcslr4zaAxZKdmNSoz3FESm5j1DhQ/Fzflb+UPP+iHet85YXrjsOtyvOJXHvnvB9BOWo5
dRaEUH9TJ4nlNNnk9XvRh6S7aeoKwRmXkB1g5zz/4WQGSFc5LOS5d56Qt+AfLJzatmhFe6oVTtVx
GE619lKw8vLaSsB/xHBFa2Ll2yKFnxmWgxJZBtTiq3KDpyJFLTOEeKdLTSF9Fp/b8l0TKqTYSmwG
21ijBqHj9jHadNwJRztwI0Fk67LiY73nH+h1joQuqqVXknn49EwaPOmhFd7h1MF+WrH/eiLKksvS
rp7a66fxDSHTKHgkHPdARJHPljOSybU1ZkWIagjJkBF3eKABfpAz1ikg492+/ztLyN25uJRG/JKr
A33ibRx1fCh3i2OcbQp/QSGy37CuvutGSC0YNeFrY9+i7fkPEv7r4Z1vcXf6I2cua6IqdFLDQC/S
yYE/6qKS5tr35lwYDAlMO+xqirm9HG1hTATNEcTy+Mh2T/xD3QQEHAZlix2DeB8wnnMMwOhXYTTZ
ZInbX4Lku4asJ/l2NQJw6vTX9uyGaJs9bjpnOBXYH+RnPiCXs+4ykmmbxdwYbu4ooZmLae9948Me
l0xoNaJB4sHTeWLgysryrN6xEdBd/IFX09DeDvgQ5lqXWXdFZ4YmTdIed5+N8nbGvboEZimXAOjQ
Dh3m1p8bh4PyqEF5gNQ60VQ4ebU9JZCFI58kLabohHlgiQt07ibHucxe0f6Vx44RSUvzBHiRw8Zn
48E0W3RxMrK7zPipS1xbMbLoAZ2n6u80fwNV9dQMNbV5h+Jb+LbmCxGG3CrA+wAOvLGyGAaiQC6l
Zp+iMWEOrgc2sppL2Yz8zZQo/xr0UNoTQF8Yl3K0QRSAibaATeu+pTa0AcptK9AmPEP1GOdyi5Dn
W2xw4yaH7sj90Rl+F+8uph7CUMsmQCuIAhAVJY5c1IkS1j3k5hM7I0tRswKmA5Hg9gj2oZqu7dUw
E2bcd9y/ia6GWAdkhzEhN50rSEvHTri/yRWo+bGuKVL+qjLRxRwGJ/bEfTRPbsQ2Fat2xwz7WPir
PoshP4/Q8eg2CPbRyjOxzsYUiv+9EK5Q8BlpXhpF98uFWlmili9AWTX8GoWhZAJXnFqBWQK4oqmz
GfP2F50h2WQ0udpLkbWeboQyH33uS50BEMCk5lhE2XPZDnm/roExVoyczowV+wYWKc/6esmKlMuX
EJujMcgASKC3LlYG27VpZToWefOkE3p6pgYehqR5DU8L26LyXBEzNWBAdq4mwoerlhqmCDI0mWUW
HzVISTmaTjUwNwnqoJG5LCSNxRaW8jpHuuAPUl7XRjdwVJOceq5msKrCz6D/IhB+vhVZmVQxrhDF
wLGJMaWzB88lf+5WGB6b1Cz4HaCzSxy7OZFA5V+KbPy1tUCpqx4jhS1wowKU51kFebd+CMwYTkLV
uv8jAaZ/KLjuAucx3yxyMcUndd9MDHybt4hp169KqFM9mcplY4PdzI4sOe8uZJdNcOYIDEFx5KUV
l4KWFjqenGsYqR7G9sKXlDPB2b/SIhj1MNfbX2HZAz9tYECrsf8GveT51NhsY73JA4ecJ3w4eXwq
YYP158ftH6ksmqIln7zZ4vA0CdWXCJ+FBR726eeDiXCtuYaLGgpZjUe8tbndmn8whEOIjkAX3jFO
qY3YJsgj3jJ8hu/TRNBXadVM+vCtTvtt3/EFuPKIKZvMewXnJDJHbQ0H96D13pojZJTMerJzJBpR
V3jbJZ1Yr3tVDWyYT/Y2BTP7k/tUbbA/irqWCgbj51P3irJmdyBkIVB/4ERY9CtfDIk06FnFI5s+
AOHtWC5e6yDzwgVofkD2djXNHBUTGZIO5tm/MyAyguuxjaA2cJ9hk3rPx9WKRZu+R5Zw423z6/rN
k9su+9ey+32T0ZkJYHbQAtrjK8FcCjmkZGhofRBG4IPSgTdRLkM8JDqd8OLg3ZtdmB0ybTN4zHoG
RQy0ncO8Vc+GmgovG3vnnLMT5dYYMrJXTuzfddn+P9M5oRr68kQQyjmoWqbkAodVsAiQHqfxv2cZ
dHl2TiwG7V/Bnfh3iRUue5VwS3B331hzhYnsC/1hn7PRp/fobj8M/SU8K2o77Msw+VkiS5qHQ6Vw
cjylcxqGY22vck1peutEJ8DEu//X3+xgNVyXjkFgZ6J9Cyd6TyQiiNVanMhrJMz+0zlZ3ypqQV0d
aSkYuOIGedytfk3rZznjnS7HMlRnIG/KPLAUCjUzUpl7s/xMpkx4Esmx+qWWssy0Qc8CX8nRWS9Q
GLvFjC/bVDhfdgTc3jIJmk30lrRZ5ah7b4xtNH/wUiHV7Jmaivs5Wu6G6zl86YTcxmQMch+O1CRY
c49eERp5h3LtajefP/Inaom6bBzXVfmApCMi2AJ7DU7HIGioHFq3QdyInuu7gGkpVcQ1ZZ+bCIML
NtDUvKEewUjbN0kb9ofdL9e/TiLTZHq/bRUx7t5j/tOEOzwlPg6PFFwxrH7wF3dbCKZkt7TNcvNM
XwINEenEc3XS4LFRdvtAgdGGcbQHWFV18TXZ17e4F6X9Qs+zLvK+4L1zXn/B0ooqo9NmoIz2jwyg
jmZ4WJqXBOnQ++Reg9nqzfhDZl6Y06Xk7vkKIOzS/33SgW6EMG/wkQXPrLnNgahGvxZ8qfsXPwF2
nXLHB1FMhwXsytLRy+9HB31wA8kJ6meNEwNAKP4wAPeCL5n5vwKuhVTkfJ5GjU2bquiu9HKbw19z
/zrLGVPhzN7vxnM0+mT1Vi5oeNKqZyw+tttCRp68/De7wmRI2vZr6Sq5Dfd1HslPwIl4q+IAwF65
oaSjSk9lPoZiGPjvQacnFht/SxKYVS85vbh8fcWvsjXnGNLIJTmbMLetlXuFDBVzOqowE3yBHfc7
JdvbeM4zCuXhvA3QwxIfm1pFaVO0xyFOIRkKwc0EFWqmD1X7m4QyVeyFpOgYRaL3EEZPEtp7SvUp
muicQwMAE5oXWelMXFeOHHQJDLOZpjgIrqrVJQdOqW/cmligpn+bJv2dnkWAc5upvXdR6aVt7yDJ
V+5Wcc2xVDNEs14NpQvRVdxPWVou6GBmvA9dPuOuxASdm/gf6IEXGOowJcSigR4MZ9qgVRa6SrW+
1bJkZEzA5lzR+ku706AfMGI6KHPZ613fGIl7pFeEhTN+6YihmrWMP2vcytEAyoQwcY/8r8Nb4FaU
tYfzIgYNKJkMd0vjQkT0//37j5/s+vKDq+klAbgrHOvKt0fn/EE+Aoj9WXqFHMO1W5AM9L/l1Zv1
Jov3hQwWSkRVrwj0GOGo5tbn4szygh/5UY6jWLPgN+mDbjkXf7FhoKeoic8cxxEFIDvU7xCQhB0R
6+/jsN6NFpLA964oWKhNWxxSKwmsbt4YCAhDUrOoh+4mZE0lQS3eqUF6BSqfu6Xi/siUh8W//wnv
iX0YyXvOBBU8AE1G/P+8F/bFWPhe3npA+mlZEhkHdvW8QzaZhAl99edobAa8IudCRiIfJrKKNpTU
wVR3EUEe/KoBhm5dyJN1BIWUClHQ3w6jwfQVoC4GKpgCgKmh5ywZmNoi2Hu/7r3UAAVVrICQDTll
xOWDw08OpKFyzC2MnjIV08tqRs/lV3r9FmbTlnYvrLQbGGqNFNYeNg9pFi/zchz+QlB+aO0b+tVl
MO9+EcpOI7rKmYwwniYLfWWviOVK2ELJDduRAgDUvouU5x6xfpCiBElzbQyV3pfq/Ca6YRTgAcsH
bfPmRxyn35w3TLs6hrH/QWeulcTxpKdVeV0JcgZSGRZGWoTmje721T8PtsMfKJ6KBU55VZ5mwVLz
+R7q+RRW5sQAq4nvW20EcLhXwbcWnvjcJFCrxGD/60qd1aMb8au/MY11j75kVZXKgU4oqhbx8vb9
J3vSMrz6h9iik41W8q/zMDt8zNacBpKpKipz9LruVFtMirBDUhxfCVyhHiQ8m04aOrTgEL2e4GfL
+VPWlFmZCams1Xbf/TFsEoNbUfKI/b3mmUHB5JePvhCBoY1dDZN/Gq1Ca6AlpauisTkQSy4NEvnN
gzKvNfawFTgUS5Ay21IsFXUzC4eOeOJhkx8oQBJ2Mlt3RkVv1YxxJ9ZhhXkh43sTugOE9mSkpSmq
15iKBGwHO3tSULkiXccjYhydZ0MhHpySFykuoXdC0YP6iTKoQlK6W0giOJwTxGqVuafZCnTr/wmS
gn8wxGFif2Fd1gDcPC53rTaSdt1wAwWr28VQt9ohxg2Alv9QH0ppnoHZ+AKUzlbbXZtHDmxbV5AE
jr8K3EzXFtta/Nlaqe7xE7RXObJVl7uz+O+DhvzJbOVGcWIJFFeWSHAnZqRJCwY86QeiX9ia4kCg
VlBAfTvbSGpCPewOJzBVLjnhyRzgwu3mYsDt/LH+wuSXIcRwqXYn2Qa/ZqR+lWRIf310VJwi9S8E
PlRiv+JHncrge2QG/9EqECAqJH6Tdmt5OeR0GJcr07WbZzz7HG3lT3mb7tzAAj+LY5yOrDfCHrg5
MMr2S7QeV0d+q5wIOmjwfwajyFKB4LsGFxmZ4zFHKiZ8GwdaYelhKuRgxeKvudIdo6rNAKrNroFb
4Xfu8FklsvO9wa66B9SADwoyYjpMEMiPMR65iGlaRJ0KoeTBgrafkwMQLT6QrQKBthvXIpMSd/jA
a7BmYJ2Oj8X2ve3/9Zf6li32+e9877DdRyZ1Vk0ammxq9k24b4mCV3vro1/qrknw5cgKC78eDu8r
HsIHktnyiuuMi63OGbHG27B3iiwwqFoaDIGjJI2BJ1fI7C6IutxOi/M1KnObr7vy3J6ljPnX9Aex
Vz99A6VUjUTHc8jndFyaiJutq/YnZejqm5APrfGYdbezY4g683dItYuobz1JCh49VGxyIAl8+1BZ
7N/4LQvDneMofXGZFZBUwXEz8iuyOZ1cFJVsqSlfk6cqzFddAJVT+J0nHJdZGKPfq6BjvBK56IrR
rs7fjyrRIZ/2UnZ9t/9uOLCjeUH/Rvu01d8/R0/Vpc1y9IubzqH3ZHUWCeIt9Ylc08ZK3Fj2MXRO
Ir1qmELldoxHxNFNFys/3Z94bG8ubEEOUhJiIoA5W5zCHvfnhpr4HNU6JBxyKEeSbjQAWakKSqJm
QZx2TOl+05ryh5YhGpmnvZDL0jZthqj0w3LRaOLhLfXGFCKn344GtjOgPaCuPLQWbYkzO2eg9vBR
r1Ob6H0d6tnqflXNrveaw9QcjlnqExZ7w8wp5JG5UgsuX2UvkEBW57riUsnzavTfiGcKMDNuGG5b
atH3ibD96Y+RGBHX86Up+fhJJYVoQKTXqYui1qB04TQO0VEzIEYcEAW9X9FHTL1O1HQR/fcVQPbJ
VS5FcKT5T0DryWiHILRVHXZwfoTNKX/84zTCrnmbfyeDq05s/jEwnGcMbu4IzA+7yRiQzXhx/8s8
CpsCX5JlbVqylC6NdmndcF556HzlzSDlKqlhyZHZMmnP3BPzLPZqyyaLEKpVbTG1vvRJQ36knKp2
HD12KWIt4ID5s8PKZZ6uJ0ehsYjZXLEV0dFAiJ1AELyMIEPn6HfC7BCzRzUswkdswrXWrJGukEoX
3+2PnLASuoKVz9CLcSqDH+Y1Y68/eRQW0qKsvo7RQHbjpF+MzkopA6ii3CDZwk4ErFGJs8Yy8wNT
fjppLjCV+QKKEim3Dd2SWtusOG2QL0QKyFN1Ded2ghi7DlvG5+MEwZr9dBUh+/L0YLoAnNpQjWKI
dHZ5SdUPRl9eWBlocgrfyvaDC9BaPfTETvrtqeQsJBWqsto8wfKUqUpgR+XPvxPp7y9v2CsGWrwR
uQc2O5Ny3DHB+ohMaMbOcVZkE1R3jZ5XgA2++DhpDtPX0c14ErjLQI9wqnyZ5X2h+8BKpw29zMqh
Y6L1Z2nlPfGqV5TyHoxPALd+z8eHQAhg2msiRAmjd2zWZmFMM/a2nFuiUFFs+fE7OxhEwhNQM/0S
mJuQRlM815L7AlNNIkJkoplpRG5GxH4v/E8mmdJjQz4wgkau8r3dl72Wq7y1mgnNYerhM+1N10CH
EFnKeaH2up8mTeekuGN3HPuhofXNV+dOqnBKAJw5xghVvuXPEfY40MpNst4Pnz3lekanTFHT1hjW
3U4VV/HMXmZPq1VkqYdWMMwE/az0+LgrEEC9YD/5wbqV+RTqH0sHY+loFozn5EdxrmFVh3CqfAu2
mRM5jb5g0/ruF2F67k0hDSoCVq59SdTyoXcTVaoUiakXba5a/VEc3PWbNCxd1BRGu6LvF23kZqDt
m92hH9wXylDVGSZla8PN1qsrF4pYz6GH2fh+yGP18etrVTTVUb/lKpUfQ2UrEzwZtBzIGm/ErIpB
Atyh07tt6grD9T8+Qh4SKEHKXGyW8T0mGyM2XMtNXTvF40ONXq5mf6Im2bsFv+ZaenCe+/9WMcsz
tF2sbr8jT9wBFpAbzQd6U0xJeQEgjGTyvS27YTOp1x40O6HV/0h2PcLu9qRXh9JmpL8Ik9BcNDfs
wyIcueYVYUpKHwEOGrKwARFIKO2ACA6wDZr/6nCy1WYJX+Hdu0wRQxsM1i+QRfYz9K90yneoPvkQ
ig6YTW+Eu+z5E1vhLJdLUqZok7lpC3N8V+N7pXA7BjvYqCDxELT5B05z+L6xFuzXvid4xFKT0F/O
aHkQq8TbCd0NIKPvc9kTIWTEZaYJAzj2GebDB1WLofF5nzMewNnPBXJd/mgB9bbqTI3FAeki+bVG
4U6KFGIdg4icJnzGGOVhhGIMRrc09C+esHXmzoupKUXfBgaW6JoXkGJ+G7MOKcyqFPXMHsJ6btyK
EGS0fK1iizMetPMlr8f4qFYX4abQ86G/TwpH7KhrwNjtSnnZXd+7e8UXX6rQWb/PZl/QwubaklBQ
b734/WPjy2I6D1W3xXNhuhmJz1chX7dQ7zQsJ3lVo7NnSqGu+/AxuZFXZfEVcoc2G+KkpMATAcpN
PvecWSTxgOImltDSJ/mNfroktsVeCVKqil4FPdu0+/soH5molzRf7mbOwsV9yuoiE2Rk29Si07YA
64/ibG+1SIdL+wfI2FmpM6W67VPxhuthrVx047P2LHZcaiR/zgGGFGMVRyFIXYESikQXpxbEtLzL
5NKOz/1GQHg9fh1e/PVaRjCv9FXTS1plrCTgb6MweO+7U8KYK72snS7wrfoe9UFVmpe9EqGH8A8Q
KdWusFopqqCFgqrf/MxgELnVSpyW2wFMQtzAeFkygaGNEqgRrIxCPgS3/JDljj8wU1UQBZLfUO/x
TCI1Grc/uHIGILBDFmoDCozvNUn2QSgcTc41H/9I0s6JsqLpA5Y8cwVt7yZF3M6SQKT8duyDGsdn
UWoBGruwhZhzANlFKG2SJBI3WMtO71rtNgFRqYtiOq06CLOn19Lob9pHIetSzZdZjsi0ZFEwSL4O
oWKvWncuLRy0s+vxQXvHBklbb+nAoq9IK4roe4wWBz/JlBwxzpWRd8fyHHfFdU+6lON0zkHBMwdG
PpueBX8nAYnQbAX2jXWBBySbXIeFGKJK0B/QMo3ocNhPxQgzV8Jkj++clcY/WtcRB1QNaHeBp5jl
9BkdO6t8aiXIj06SKOS53AuFZkoQF3N5GOUBTPoKZjiouVPr4s2q1coLu8apg/fVd/ge35caeo+f
2cl/WHxaoOG9nT5UP2UjYx0K2ntrazwpFsOm2uEyvT1JP3vUdjG0A0QSxvOEK+hJlQwlsgs0vqef
v3S+jIuAkTSgnamThECBxQED6hXVvhViUo/wjcAN6YpTA85llU6xFOf23ExSvgtXPDBERBjpRGLv
KyQDnXaU6p1TSIQ9pLKxmFq2xA3r20yTy8gXQZ94O3auFZAZFC3H/T2j8l745C54d183uvDJEW2P
hPRKjDKlpwKUOeYGqgviwycCEwcSGGpO658Z06tsNnKLjdldZRjxnJy29SZcWPbp1Rie670LbHeN
v6n4WZcl4VE+85ZRaN2q1NvjkJyRQURpz0ld/zl1o0YGxsgLMN1qv7RsXWicO07xCa0JFU5zz5sL
rA7ZaqreDUfB9pMplDAYEa4TFfui+Em+jyewC5SZEUfuM0L9/4W3Htmd5Qkygbn1KC53rZwh6jkg
bFLyAxYU1E5L6Hjvlti6xLw9HPMiQxzyLEOMjgK1AYLgSKkoN8qWvKG9DpSl9ELV1gK7tzd5Fdof
b3RQglJGowlX9qLlDfzwtQzTooktwlInpf+uhjwOaXktDQYbYwrdRjKsGfHsGc0/JIMgRaGiCeBF
c6kqgnDdBIDa20If/FovvfZKfbUA3/L3pVVrZJfhbuYq4WwVJAM8pX7zs07gpLFYVGLMOKvy/PYR
mmmzJk1IGNefcCHuqV5welQM9AsvVR8PR/TNKBUkf4yBofb3qfsYKQ7+S8wmmwNgsNdTd7Ka5CjY
tQ1cP80dZlf8lsndZd4t0vbdL9fd4EZ7ch+476B+LKjGiiOlolxvpbHIYGneTTTj9P21A1r9Zf14
cC7ATzsuzdBzQRbW38qWHHDShE8ZlkmwBFvLjYoeyxgwH+GWTRlKqy1eO1rh8rHQobN3+go8ikLd
PXxhRSoztmend3XDN1+n44YO1NhYdZXQdrx3E5BaIbErYgtImHwViKZbzkbokTkjcMZ4xRTw3iir
UA5BmZv65qyIJ3Npd8lGlVzBLDMkuRf2nw1RqhXtWf72ZAtxWQ0n/Z5ZhupqlDV00huCqyiJP19X
CkKleJlpX8w1YYgLya8nlQlhf0o9FFadbepAbIsf40ldAEp/iZ9WYU7h8brsdTpqvoklJYAHD2e7
8aBkgr8aG4nXNKUJZdiB+Vc9hUZo1s8LNeOs8zkxEdRgJFDX3ED9xgpOeON4uL3ZSZi82MvNTSg8
EUj/gwgvICFdSxaetUf8zq7J94XtIEUVHRhvF35UCNSKNlux2sjBcTzcDzy7Y0ZKtiNNCpE+vmhj
3le5h06QgJa2xJmqzlOEvOA3tv+OIeXGgKSJz06APTnS28LoDvJmaOWXPXIgtrPPgFNg82OlZdXC
+MixE5aU2xesjiejv0fHQjyZWYfmmS5kT5y4EAecrMfFuQYVqHb063oLSt4cSRlARY6TACdWhOKe
BKjLbEGI0o+LflbufTMkdx7T4gzGWg04XsF5o5marhhWPiHC1rAr+nOiR2OG9t0OrluH+HMKHcMF
yhkSJbY2B/0LbP+Qdt34wUmY97Yt+ob5GWeBah3eVjLUHEXwX72GKeii90zvQzRDgPiaDPg7rJOj
J97g1EpGXhdK16h8I+qAiSxuCDQ1hFVZosz0GMLbOhnSOGFP8JgoIdLuACLHKDPC6UXqhM4zCXzj
r98LnTsgETiOKbYlWpQ81NJqTV8Enq1JWLE83mkPEzpmewX8FUyGN38JjlDNjlyTp/5ugtImcmWk
wtxg3KSe5fMDT2X0DdQwpU8cf1Rqo+aC99IPTUosf0YRqJQhwJzKpY+Wc/YhoiIOuG6up5bbuJgT
9WSJ2rbpW9/f+t2NAESWvRj9GX+PHRsdU4geYsv3oN3IsW2sPHV2anXhCiQeDvB3uUKTknXQn0qS
ogfTf16osRdnFdBUt54JgpFpqo2ecrJWFoU0nZbb8dOvp/VH7tbpTXxSu70wP7uKrlYBU2nnG5IU
+Co+Fn3IOwwIc+zKWjmgdBr3OFWOgsFOcr9wMOdNJLP8OzzMTApV+2Me5LnpEKgbYVg58rekGZrq
cWP4hW58UKzBZ90zkLumxt8PuVBgTuKVqPfSaA/Snx15zJza0DJRf/0wg+JXQquPo37KWFKU1Yxw
Z/XN6ElXt4r3Ddv7HPELfhCX80kQLxg7UvvHS5qf1I4spkw3dL+62Fr75Q3uYhWdwjt9IFqG2tre
ibW+zZLy45aimSdh7w4XDJPsLVI5zgAzPYDF5GuxvsAct6x0e/SROi4/WANL8P2Bi1BOELJMBkzD
ZPYfvI2nFk2/NU9m6tV4CJFzIjb6lF0LKg3plj/Q6dPG8xadDIKXEJFKc0ob9XqiyZ7+Gaur24P7
wCAtDT7xMj19DxESORpzjQtOOy6ZiAwrFXApi0NJTC33VCHqrpixS0LPd4k1ldl8xdbHU63otOoh
XVzCfeOnHMhh6OVUplQ0rpy037pxuT6o6KA6Yn+9c+DEiBsblKri8E1Y8nZ+5zfVR0JUKvTM2+5c
oZeNmBR7s33XpoY+r9k1CopCQCiwbRHmrPLEMRrLNGTTMZxVA0cU2yX9kwKRE/At5/g+xUl/IoaC
s6ZKZfDqVOlq3wBoyO0XDH1JrcDTrWa9FNjgym4LZLU1zcuXTbajZ/izu8K1i3PEAAra/2TI7Ws5
PYGHBQ9c+jXVGhC0pDwSz/e8OXFIPYOXuZy4eOTE4iWvv82EpT/8Txi0ylZi2kvZm3Swn4/Dx/Df
ZnvJGm/4FQfF+IaCHlH15kEz3u9ZAyt1TMtftZEXvwG8xRF+yEX7H2gvqFCpyoEye7yqxeLrilLp
wuyXVKrIFdhbFH7UFypb9TkYLyAv8ymYWyrLzBuMMbIAQUSBM4JectQpkBcND3lM5Skrct3k2rrc
NufvnH+mDWfK1YvhjFsNT8WEXIxElnpTiJjrC0dCgEo2jMXoTnJq1efCmLvYbcBcDs+BRxliVNNw
nCxKoSWxwQIeWWAVeGSBC3uv7pLPNtA7MHb0/b++qBY5ZsViuFF4ZeVyzlnR91Yq18nKRTO/LJB7
DPVO4ppM/mKQvv0N+uILjfYHTXpI4SSFwd9C61HdWy4EOPjbf/0KrX590RubB3Jlc2GUsQLvYGHe
A0jrJdPPxMJaAfT7Bi7rOlbLMIMGJ4RCRYDSxNN5kyz4kk2BMflsbzCkcEbyoPjAcu9CdzBk51dB
ogw3KDcBZ1wlpYnhfPV0e3Pw8to5jYmvQ/cpW562SkSfb6iuYH3E6dKZo3NMXTlNPVlDgWgW3v03
TfJn2uPL7hQpr/iJCTd8/rIyklbElWd0yolgfcY3Z4bP9gnRTSxzKx/U5wBNSFgC/PiiCCQzQEA1
gcQHdfWOkKrfT3aUqKNSL4CLXfvearNiCw9rcX42kassGs7rWgksBq0rq+7KIDsqUU+RyCe863od
CZRv3op+U5sGnboQZ6rKtogLKFdUP/u670rlyuMWzi5pxk1rxkFKGVuQXRCz2X/Lfs7L29bEPRXm
Wf1f6/woIlPjyO5y+b1ppMFIM07TZS5rP6E4CTOvEgt9S2tAdpiBQpFHPQNUqLYxaIAJ5sm4qfhe
SOggicT9WwaZgeH0l/pS7E9KqioIiJAoacOTWi8RvZzJzawcZ9S8uNfYfGkWpX8NFKYRoTXzVXhw
CR5gjjJeAp/1IAqNn0h4hONK4u4W+b58skerYw+q9QDX4vTgOCOLANqH0n2lN0F6io0lpvRg4/kx
8BkPLWl1IMIJD3iFIbjZIPTEsRJzbkdQgULBmiaoQAM26OBTZC57H7lSTmYLZybR251gpyMOhEbf
h7dU/oBGBx/FbOPCWrR6PWkn8OzDHbBzF3rVGyypxJwISzNkI2UMqRsGPWhdNTS3QEh8oRbiGm/m
bTWapd2KzMzxAhgGkmvdJo1HTEwHL5hdVNNG2PKe0RovMM6eJhbp793BfRvvsGBXnaoyVZJD2kor
toUsTzVteNMSr6nTVaMN7F6wMS1smpLxjlcyFH8wXQnNeKKCeuWU4DJYTPYG8/TwtxLLngCo0RQl
rBbdcdubAfD44O9/YMGT/AX1grdrQjZDmDOjRDpJvb855VWE8zhkmoQlXeMwCGVdukYPKInasJlV
BEhgFUIqNZqk46yL3OKJHamZnMv5asePvn+L0nW1Su2j/ACUCBwGP/0npGKLhNpR7WLgZ22Lu2f0
8TArTq7guJK3e431y9dzg6Ay0AJe8xGRQDXP1ySOnpCFv5/SA6MVVnVRgGnN85FnY2cdygxbK1UI
s3sUCnNNh+vtbbH4ALWqdaIRS0h1jh6jNwdigTXjjc7qIQIevFlHQLMhaid7QOnjDyIIFxtGO34p
2nd7q2eJjGfhsQpVeV6lITcbjdzftnXY7nlpKuMe8bJvVuI8Wdk1kQefd5pWrDNdHSxf71JFOgIG
l39gDHhyIoHR7EuUDbHM8/NdzHV1ipjPNBM59k04A8V27o/JLGQYXd97UyGINkgMRv5nA15DvjgW
0V5gSaA3IeOl7FSBzX9qbQsVa/06TiNQCK/9S71lY+Xc/TP4xpS4MDOZnTr4nFYtCnCMF05cetW3
5ejs+uHpAvi3/X1Az6s7xsfEN3nkNaPZ7H+cUQ/yUt6CMBsIUkVKCtQwvGLI6cWPeu19WhwGBP3+
Jh/gEKM2PF9pTtPcx2LjTu5WSRZDemF2Uqhu39e5MbNzAmbDphdODXcjVM0OiVXJklIo8qqWFPyb
K9npMNaflExAv+BhOlIO9K8263dgkAXlrKUvFd0M4Zb7xH8vUZXNaubZqbwJ+ujoKkvwPtwRhp+v
cYUUwDLTTbjqrZbayJJRZa7MF5fDmCItgqwa2joOC6Jv0Y33/IyHPRpfLquFOR84vTxWOW2entrD
/fVoTxoCSqxyhbMjXDfmqpZv6mf8Ukiy5LmXxtHZfCZlnDr4Qf8q5dMd8JNnuLt2+ooTn0oB1y4e
lvVuSElMut4qXmxAck82hbhUNtNqCh4qlSlM1/0vBW3SKSdD0S9IWv0rv/AxzgeZ5W9/ZYV2013v
wUh4nvdkMSi4UIXUrJeeCH5tv7d58RcZLkfaIVAzkgc4LGP+GHQGyZftkBKyYrgOtif6/8GEbAiL
I/B6pZr3FAmilYA6XGg9IxVXykjckutcGNmkZYtIKlttqH0wV7AKwKwkoSy1yYshdpFPN8kSzLtU
Tlt4Ix+KKmwVaR1uNyHOyleoJRS4cZfZ7isMWPl8n2cjlJCmLxjiZf+7p9s1O7fLUdYNpEIDpyJ+
PVU+ndOLvSsmTffioGfFJ+goElU1yUKXn8w3vD9qqk2DO9iLfFHa1qFMKvN0Z6Ii7f+JeFucuNZm
UeOVidvUKuYvntYFturDK7qJH1LTtcVplmMKFvG6x7AAUZae/6o5jOO0LohqozP/DkGUZQfrBOVH
2Hc3r4uirtJvt2S9D+jKB8EgKZOqcz/7jM0sEFSbQd4QIvGt75hxOuhFAGkLvP06U7ZtYpFj5Gk6
mJRAr8HBF7IfslwRh6qXLLw+7uNOyoBF8SdOK/TW3dgTcchMXlewnealfPSKNwIR87w81YB9Xz83
MZovwLGmO+LfJR0nRu0PDjF7nOZIZeIuzXIc/hAQ7QtsgSxDz0uxPOIawOC6MPFH6ofUpsxN+5r3
uODszjyVDVqySnPhHvEmR+61pFtkSnSssxr9tIFo9DioE/NK7HcRRVdibxHUxe4P6w6DMXmg2Ful
bhUO0v/bBDDPZ/h6QdM7veJHVfFA15xezg2pXWceDNa/duXZL6+m76bRWgxu7nphTEgLjTpsM6l5
P1rxF0URdHV5tniwoLx/hO85C5MCeQ2mStUaHezhbwrm6NIbz8lo43atv8CohOFcEevNKlS4EHFy
16EjGTykh7EH8EG9/4uHB34IUzOP5/QorMQFNqwtmu3sIsxhlDyuGFgXSoSKJ4/x4dIBBDCd+DCF
2/bXB/e9g/eUE4iAIX8tnkla1pdtWHFRsJ4GTtSF7ROA9kBarG+zitRnsbqKJsvnOTVCQllgbP+G
wncMMjNJBqZiUyMvnGwTqIcijIYh2Em0aOjtBkKE6iuE+mXTUnChUjAhMhxV16KIWVOtnulcwuo1
CZdg4FTI9EWk4DcXKu9YphbZ/dqZ7EqOD3PYxHI2b766mytnJy3IBORWK60YK5Q3bgts2jmMmbZc
P7rqKCAudHyidZ1jpOWy2VygXaqLUBkCvWQN3bZAJ3CfQ7A7EcYUsjGIAEYNvlEBT8Dm0lJWG47c
8UXKvyUp/2XDa8BcKCykIhdvTKGVcq7V9ZlCAZyyXRnArV/7KoKIjYrs8GH7loZF7dT92mbdAwYW
eh85YuaZAIoQnQzlURsgL+WOvvG4mj6BeuoevJjSyg+CTXKi+QZJ9ZQ//YxaPvdA0wi5z1ekpBZK
ACMgNwuqVZ7xvQO+WqZ+N/eJtzFijIukQLxCahkalAsnAXSHzYHXAR+qwUxd+l40JYyw1B6zG86I
AUpRzP6t5yWURE9q5DrV88wBcgJcF6APp+KZrmFFDMCiEgKk2IwQP4BhdaYCRLwjL9/KHXUJ8vR1
HGoQiGfsC3jv0bfsvi09nPLLh0pDv02lvrcPAERvPY7XWH+mIEilkHso3i/1sBCZshPyQDj3+VgA
sh58g+WjexAvhqVUSwJLJaQiZr9o12/er9KtIhCUMQ41TMaV7Nq43xWC0c9SlgM23lf3xV+Y9L7e
WLSa8lxJuYy8A9JCxktoIIqs2LyWpogeJEVxd32PDVhT1ivqene3onZg0Jd8aDXUUOqLmyOhl7VV
S6vL2g5+pDlNNvIS0E7YvxC4QpisSEEmBnRE3EE7OFF9ds8tmdp1PuhGhag3UINRoBv1sRRPHGWj
driQ5AG1xxzc6JbGdMBEWuoGHwKE/p8LA3r/NkQzkP0Q/NPrMUlI4rru7olbzYJf/zKcbRucb00a
kgI8lyA7HyDhZ0RyEaOIlGxqVzjhbRKAugZQ3qMeO+09A2vEV6JKcz1i+iNWO+nAeNPf88IXQzD8
y8LXea5KUMYQ9OjBtBlBSsieZeXPuoeZ9EjVhPMn9z2f1DV7WWwIF3QVK7Xhob4GcsH+DLElBNv6
hMujYRZtxEG6rPPrDUm554cYl4bSwbCkaqp00CB7WH90wI3VpWN5SRJdmBtfqtHf3Il63LlVRZEO
uBMZlfBxosAbHdCkNbLrVkqBUmdMprSs7cIDvW1+0fV/Kn3LPouiqjj9BjoXMrE9Vr2DY8pV/DEp
rEdsOyRkTessEoPsDfsovpt5Ls7gdsNnjRDp0gNeO+rASCQ+j48uhkfymnYFf58UBZfyLCPf78oD
xwKFvckdNMAO0JG4tVdSDvi/H/UzFzeUuY/S4vitcDwLv8V8PK8VcxgJc04M5Ya7U6UB7WO2+Bkz
ProfbA+8USRF9tZKqkpNxqckGQNTllJTfoh0c7x9kC6q4TrbHj8OSpPOWUQtlR3StXS/ZMYP/PUn
z9TG53NLM+d5J7wD1E4Z1zPNDjmobgXYXzK0BpDP8U51j0bVx2X3Qm/qcwtg5OzOPR3iCv/q4MgC
hpU7oUn08Xp4D4JqqsaWHxHRkYYmI382dXjttkA473JO4zHaMFZVO83kFpshDXfFE3thhP9P5vj+
vVReTXWXthudT0ROImfdkoPY8dlvLgUrLO+jZnKO0AsN3CeU7dP8gU8fb+M9llWWT7y+JHRhZI6Q
XTqEZyamkuEKmEplupNJgnYMI8kj5MdlJCNJMqhFReCMx2JaKZOU2gN6GUjZjSAqpBCyP2mV2goe
Fb8zY9ng2FxVhCFJjgxIEtjO+r8XKZJPvz/wdyFqYHpPwJQDpCW8RHKJmfyDFDozzwJ124+nUFXd
0c8No2Nof1nkwIS6RF/hHaIGqaaMzivruCDx3/vii8ZDhiQubCt59wJZd44XXIwAkmrHon/0T1Ek
gIa9K6uu++Ofvy4JFDmk5/1cNy1fSbPIi+7AnhWdHTyl6LrcbBz4ztDCHLUmivxHabTL+7YA20AR
Q1Afx/JCg2hMVP4iErYJnNoqNLQN5ruy5/cbihLoiGp7XSuY1W4rnhwPHg+xb6RoPUVhET/2HlJ/
c/N9BIkp4MC6Wr9LrSqVbvBo43ZToB119bGzqeeutB4Y3H08ZKq3s96zgxT7zonBRRi7WWaLcrkM
GzQIpgvPtjQHbGY4uVHKv8+SjDbCzQHPNGSgHxNav72E4GsMTccjfmWjC369KYffbZpP+b6+90U0
kVMH5IT2LCUrSIK9sVIaxRJ+F73ZJnol1jPJkUyMnA39wnUrEbvl/4QMtTy6/QTuW+Qx33KT4Avh
Q59BpLQqRezKGTwHRrxkB+1CF2WKwWdDhAp0uu1JMmVrn1J82a0SPwsgyfNYg2H5oILff35UqF69
moX+v7KO4ekSmVCYrhPjgHm+ObWZ1T3ZKhcW1LZEtAeZHHkzVlSXLMnfmW72VxenvkPAXN6pdI53
/fA/UJBv4Pi+cybHj3ECtoWknZrTRJsBM6uHtcLD6egd/Pn5E/BfJ3uIIvPOXYHTmdkXmPK0Jkmx
biiSTEsegAy7nFpez3BYEkNvqG2h7A/WugmGsU0Fxu5oTP5ByGP9vDMZqvJP0pHoYnACRR8Sx1hE
X3Nz6QcLEJghdhSkeXlrgc7jPr1SViQBnk9Qzz980Pgoh/WhNuX+FFap6lxf6Uzqb6ISJefVszvi
Jj8FlNZ4TGJqDiZEQ2yaRYNGq+QhtbPcjOs7T3l2NA0YU4fXw/A+3uuD+c7yODc8lZKBg0ecnJlO
1pLb4VDtAUJK/s88C89EMfQ/ig/cWtD/YmcXjJt8m0NmyEYS6xoSDc1TdgR5J4Mr2xpBy0lZ/G84
aL7tXtrzqeAzops2MGiv+hZJLhcD7MXdMrfQ5JfGG9Q6rtQaXqcby9hi55ZsWgbfs32zOdKyqU0H
l4U+XVE+rSbrVoUXLPkqW//aWezRswqSrk8mOPtWUHnL7NXCFrLnEn8BeD0V9F52a/6ub7MQrHHV
lZk/H5f6rRwZM9OgUIrxg+dkBG+UW6kfAmCS4+TlzGxskklguI5suGFIVCOnda1JOPBGKwOM1lXO
SsiHnpxlkNHjXDwcnjyJF6IzKUh4rfeEhwfNd9OefMKX/XFQZXxO5vfs44bwgU65/JNURdYHvSZS
CaACzpNaPh4VF3XKyStdPmVytpVUfosZs3eOPaAx/TSCWkiTOOmi94vwTQVUdVSUzWxd+gy+Mv0y
kdw/KbyWv5Uvn0xin/iOk6rAwniDB94549iJiY/LeiR63bggKGSo02v3WvG0E2fr4bzuspy9HPx/
MOviiJQ1G5fUWtFWsUDDLeM9SKDAY44RsZMqeTn2zF1Vz+tawzoRm36ZZoVUHDTnne0x/WUTZYE5
VUCVpmPWfovRCb6AQSUsMrRCqbdg/33TPMYnggrK8sEcfbfO0r8tdWYwMytck8Z4Qk8mSb7j2Xem
TNeh905GlXhJsgwavMjvFFMCCP1zAQ7z0c0Ygk2cTa9v+hrudeO2TbpHpVyFv1zRnYA+aW4iL7k6
q7xkNKFuQPYqkKD7IJO7IfgQLREUoEsJGzo+/M7VvyEN0S5Cl9PX5PSnMjvpxMIePNacfzekRXMK
lnwq06dqvPUR01kNkNo6PDQDXhQzyOGYWKjjB8lOjyLIRn6vOTKlqvt3mIYq3UUHgF8Q1Kky6jIu
tKBtZN2MrSEojMjGAORT8b80U1uCGGLdt2+1mujjJ3SzcVXCWDVGHeaFN9GrTY0379MPGGZhDeA4
pCwcvG6VYzezlSnaVZvPsvOk+56c08oFLKkK2a8aJzo2LuiYs7o5ku4WZ+tjwElPc17vkzqRCo2x
/qGIXkUnB6jRlb1IhZObmwYxw+hv4zRkcnvXjLTvH3unCOla4qxaTpOL2pGBXkhadGkF4VsRWD5t
ac4Vo1PCUyZ13wkgEWbouxgW+1jqRdkHnIABYgcd6F8Zcmgr1WthioPcS6T7E7NogooUlkpimaAc
kKoyCIRhT3oEnVu8qFdzqXXX9xRu/MigPa4iNadQjvO2hQwSfwb/q556xRCoy2d04mJrQWYLhH/e
mXlVF4GmfQC8moLNTL12idlymKv36HQ/CH1O6CsuCpDpjruS/auR3hRmcOQCExG3UdeBuyGrR7k1
YKreZ1fl+rngVMZsNnMO8CLK2cbgeG1PwOpfKerH0BxlU4jePJnf4XfqYfl2IzALuUX4nqcSQqrO
U4ElGm5YcVofheGesQgmwvuDXN1KwYlF0WsyhNXoXKxxTUexgnSKG8Lk81VIY2sbkQSWpAgxpUm9
gOzVQwnDDka480c6H3/q2S7oGaffLx0jkwkVYlXeURn00pzB7QXMRLSedEjdIkPP402CcIbDX4fF
pdidfZr7oqJuGIMm924pf7rMn60iB44O0ja21jqAGyZNru8Zl12Co1SmqPRv6fNUff/QxK63YueH
T4iwPI93N0/AfzxFvBKLEmQlTOaROu5bdVkJBV3JqbYEF0YvdJXrItbPx5PEUEi5tPqwB901ZgST
nHSNJDMBfdF/OhJOyB6QtKPi39WsqanvnyZfbUCf/vPhj4ns/ym5enPZPji9BNQ7bPnWIjyke5F5
v7xORNvkQ5XD2+SBvnxNuDDooXw9ubKciP+F26w8moqroHZ8Z7+zMb3gkw0RJzjrRFaSW9Q9ts5H
xzmVvAY+vCksnnZB2mQXwOKc8iEuFRyoJxLwXC3YhBh0T8KBhcTyM03rGLhEPDZ+YeqERi7U6sTa
+MNCuOwgbNK0qbkvddUQkBDypcXEaMCAMgNF9UGfzBYMXt+D3jc0i+pulPatCqXlFGdVSpZ/on/j
eGToYqhN2ZgmxMSBl+/4NO8/E6jXrb9H8PU+yf4y7H1HxAtMikg1pQJcZwiod7aXhp+xW2gtR6Ym
L8PHS5qS2QvUwtZD4/N5G22tI1nY7ijXzwOLCPo2ujLivHYUy05ns2p/NE1ae2XViiM0sE36QzoA
qt4ME3BK9b6Iz4dKpFJIFh3xIl1LYIM0yKL1xdhR9/jhtY+ZWcgMAXaRfKADWTl61eiAyHLbDLUr
VLIrbpdKB9s79poTSvHd8OgXPZcsUeYXKZkLa4O1E9467N16FD9CKryZB8zd3NYaWw6BA6mQP08J
PbnvNN+0MrZllDahJiV1KFcoPdroI1VR4X0pS9Gv98l/OcrycZhtXMu5TB/jamjXK44RZjGQljZJ
5r4YivV2DexFOhjDKop/udUnVX0bZj0XAxZ8qHuXWmTe7OHfalhYqe1oooult1s9z26eoJ9L3URu
YlKXthLN9bKmqD+/aMQ761oz8+72iHdlfXoMtNfeWegiP7f7kTxrPwt0lVOa1BEpvqronBU2ItR1
cJOQaN1A4hHO/yMPpR6GD9dioPyX/+xqH0ALDMnso3CwhE47TeZIy+9H2XmQhYBEbbuTwkIXEwCq
gQ1dow4oGevMlrOOrPBDmAavTpkAC1OBmw8TPZ9WPdeiVsoN3GKCgN1XS386TrNrq1JIYQzSgNZU
MAKN42xktdZ18gPIN4VMjzzsp6Aku0+VOyqRQld33stf9dGby4+1Wd8x9LieaYhudho7YyZ5C/mH
vxAw3i5jx7jPmEvbGtsFbO+YBOCNE48dk+xeBQqKnab4BlqEG5gDDe9oeyoDkLXXzusIL1Q1K3MV
Q5eEIIz3VWFzgkBuA+8rA/0Cl9mKAw21zsaHCsG42m2FNSKEtQxvncJJ+XF2Cfp9HILuOfes67Rx
108wwY7xb0SnNJH6+xIPd+8u/rUuPjXBDDJOebOMQ042bXGtbOkoBWoyzftLgiN5K/68JJ7DGwpJ
1C/9Q2SGq+NKwyDzqeps5J1EOnIdhd/saFAhj8SHxp8PS1PkLZmeDgnysQ06MHPrASrFjzQW+c5u
kWeakuvoR47JNMLRYs/uf0Pcv95lHMQbGRCtyehVzorgZk5F4vwua0sdxR0Xv+xctX1GYbAnOhZe
V+A65i/ZWdDXlLqcuZnXiHORraS/MFKrU6we943rb88nv+K+FlOr8JLg78CqXNTWdmxo/SNeVCxF
pD9daGwgkCq6o1UuL5F0p2mQAZ/zBYm6j8Z/ZPWDVDyPnNhvwZ4YiTRCpObRCo+k47U86NKy4hGR
3Uu56DVvElFfJuMvN65emM4ToXXWDBQjcT9/P8DIn9MY852dlZZtE0DhXibuCQv7t43QFB+y8oyJ
O62yBZLqyFnnMOJ1h494gsYsm2o3JMhDZbmeJ5+Kg5E6w7resgtHLBUVrbZNSUrxuThmVt7QZgdP
hb8EhvSfn+Q9eZRRJblq1YOX/xli/C1Xsi5eYrDMnwVxSP8INCe3bGiZmLmCu+OMKD14uxJAV0OE
C6jZHDrqwXtmlm6lb1yGlXHhbXF1gv7WJ444bRVVndFrlr1AdCZ7AX7ECa10YlzO6K4PSuG9c3vI
0ZPuagBm3waMFOO7isII3uP8WSCS++/SuWIv82ZSucZGsu358pXEm9qpceRyuUSY0diHhPm9p4AK
8K2bkJYcMDgHWY2vIBrJXzSk55eeWN7fVjkTzOIrbINB6mk8W5jRQh0NHmOD7cE3LIwKDmiVZf9N
FMst6R1lrzff5SCf+yk7UUs3P9sIrRSJjMv1g9QnlAhcf2C3KcVODbgE8vZ6SlnPma+EM+FMYarY
c6L20D3FcAMz8HjRV/90ij5QmF+jt+jyG3m11fINoJ+lCBzoqYcjxnLrTCYM3Kxdw6soNywo7Y7G
Ar/Og7/OwYbAyC/DEXb2jjCzgetJVQdsXIILfZAAd1tWXZHVGYm2+JWfRTfvOmSDK9BAO0xdw1+p
uQ/kahiarXp4rjF01t7F8KmxVrrY6z/Yns5I5DyWAfKeUK0UyfQHHso3C3qVokQ9jssBcp4RIQqk
J2DOJTKBHGpzVGDJeQeCqrMEPSsswwIF5gQnVtTMX/B5CR39et8etQCgYkMX7nOflbNtaFUd8N3V
c6wMWMAgxvu+5Oa0eVct3AyJo1WWodt/HYh5FaAlta6Tu5GuJlTkcwCD2i0vIbmyEkWe/JughCg0
i8qVuXn2hOZLBKHXHF2duuWKEbfgnlhKU4W4P6gCCufxVQGH1IDn6yzf7WyQzvlafiDrbjkAdU4f
PqDw/3XTV3djh+IAAUQqR2NgvFh0TOIS3UzuuI8oSpLq5WtB61p6n/XA3SFd9d802cvcOCVJj0YP
Rec3C+E9kNlXlfSgvwtRTxIgG7mQHkIE5hjjPoHQmRu7SS9DZoTYU9qlv7/eV5YFI1j11YuUveMF
02eNMQRWQiDlRMBvOSvtHmL18NEr3ESK8UOW9GEongZ40clBfVQvs2vsuMH0rRX6fo/KgyKJ9KXV
PBmjGTxxonEK5xiRPxqzrm4dRQwOfkQNbI9IS8Q3wqBrzfOUPtZZozuPx+uqdcKhQy2ZUVqO6tOD
PXpcLT+QI/g453h98qiDD6tLNP4m9vV1ISBxLCvhqMAekE6PWakMsSn0FAwRqYIPrOrgpCbXS6OW
vT8DejuLb1UroEH1GTYAogCQsfkpnSIQwbnyf9z7/GgF6tbG09dzMnjKEXi6ueE5lxZmoCBTIEvf
3k2ZnjP4wZKKBBrsOPtMAxytryY7QnzIZhpsL8bX8/rSgIY7DaCdsVhdDjEj9vL+P/cr4Rqls+em
uZRBkaOuuD4frdiQ8rYXfg3/GzzVYPZFVW3iiAc3MzVDSBS+j3tfVZhHjNGUnKXwH2NlepxPKGud
F0pDtA3TfccOMGHdC6np6OERHHVqUS7sLRzPEz/qRLlDqF6DZbMcuUtHHnd1fupuzhne4Fft3DTX
RGwlDVdy55kdK4F0yf+fDNdp+EXgMF1qAP4MtPJ+3pVEbxebZtNwHHPkuzlrPTltELGr8UQej0rt
UBVv8tCFlOOu6va81p+AHL6a1rJDjSbChT94yFgE60GA8FjuazHNMEn3ir72Wdnpuy64ftgjibAD
CH52m40fPGL/Mc9Xh7BFjwYVLtMRPQZstlZlbhrq26//3/Njoh+/rOFHPFs7Vq/5LP02SR+IZx1V
uXIzYmx3z/X3CkIkdsyaDZ24AQfQ0CymNsCE1oa5nr4czFtP/+C63yY2i7T1GAZnx0+TpF0pGghI
tbuk61w8jA/1aayIm3MMIr833F0L+0YhFVToFWqzu1C3PRiHlX9iO9BNo6qsKNYEGW9JcaP/yu7k
MXcNHjGm7dgTLLzKH8Jlx0L/+UYc8+rwxvFeXoYmOtTv8E7IZW7oWjIZV+2ToKMHhmeLhJU4xh5N
TWFSrLVavk4MbuNdSV6OVIAsgouvRkTh51FTAWSZ5r41DOpo+yU4bXw8PM4Jc4hJrRsRC7FxRRCG
V4DfNalyZ6pOa636tZhnmfy1ZMta2FKid3Fc97Dkp5kKkTExFICV1IB/khUO/HqCUAUY1kNi82kt
0EaJloTC49tQ03LXz35d+efgbd5Yz/s68CDSh/sbGQbkRUxFZInCN5Rk/kqqMA+EXB9y+xxKWgDD
/DX/B+Xq0aafG+IV3tGzW70CUN4rcJDGsxQICS5JRO/iqMAYONYJ3oKJOOUu0zEdeAdXxCSpfvvZ
p4EwHrzECL7K11Do1b7ol60i3ECemERfCiXV5atVlDwstMHk6cXk9Ns6NdBW6+7dYOZj89+A3FCr
HceK0wIsd6F9qjxeuHjs1yvzC/fgGKde/URP+DYrpShuNAHabKy4wUEo+9+0pC5L3fKJfYieg4lT
+5kfwkKMKlU7C+awK3fBEJjjyAKenYbqrukCCWxPeb5ER1GuFGy6aJ7bEKWskL/STJIswLOjXqrE
SKmitPejCZw1WaW+il930hHAraJhX0ZsMH8ClXGeLHbS8r7pebY5Eg6jW7Cxtk9oAWLMaeCN+1Z8
kioDjTnxgl2dOEOTbHdrDGGYcQDJDSmn4dTk6GxBwRMFuQOGgOXTcMmDN6KY3f3QE+t8NA+L8hV2
Py/eVDqPB5P01dK/flj0JRYYrpiKnBGtGAzzIyIkjrOxvfoW2Z+jt8lyl9OypPmg6AqMPYhhfTo8
YzKS/VlUq7ljDNbsKdeRGAjj5kGxrBCoYKRHRHHJlb9gadHwl9T61oaavOk6nddNq8TDLjgqQBgU
ypY/Y93982ZLhFJ/CeRJH0cicACVB6QVGHcDPDXNKYyPh+7VP8mUIyvGy2XecT4ZVgASThpVgSeP
AFUMiVw/FEAUgWkE/5sllblpT8zrKwQYwZJ4scM/PI6Al39fqKy1omNQqB9aycRVHqwsy8Hu5lp3
g563yStbJzC7PBA4SLOcIiG6unhuo3IvQJi3KRfQ/SL6doN18622X9Zm42lO03C7+BtWHBUEltBw
TmnY4zElcW8VaFocFxaXeDLcX08FAstxY6IviBZIhyEDssr+yWmNtekKFKd3mLoKhw5mPtkeaVhG
kdhWitXMgXnd/ULrFOUSjOunhKOLVV458ZI/0LRqPxclHTlu8YyznelhNaEsAK0MhRHPM151ZTfp
k2ieW7HD0aFM4fCOkY3hTWMLon70zatnUB4v/FK1xUjgPOaf7ODw0rja0e0QfwcSKQUQGm4fyfHa
ql1B+eaC47McqngBKdXB3YIGWpaK9zDWxYNdXkgzVLZDEcf7huO5KwdVSdUIq357OdyNzqFSeEoA
BJgBmupasQvU30/x6icNC1u/msHJCLCVNVotcEfwpLtZDewz0GOrfmKyu5Uuhai8dA0kwPJPyboM
SEopn18J60RmBPQFYqh8Kmjjg/g0vMJebuD/CDX/bx4Jl+piRyVmNgzc5PgGQWmoeIF2H8CrvkzO
ldTLDlfjlG9l13PsKVKBVrYTy3vsQF/rA0jdeXdRGipdMyrCCzei5c4Qy4N6MOoIW1u+xf8MzamW
I6WU9/kWbhYuZer79brxAkepwCelS5ke0qeqH9KPnhX/L3j6PfG8DA+UNiqG6I8DlNfkJKC+Fl41
IVaKYPmEmwEkzG02KnGlSHr3A9Dkl7vSyB/Gjg9qq2tGzyUblqsS45KvDE/mgY0MOva8JI8t1XXz
iW0ueSHxTJi6lCcPNLiL3Rib7Zgr9MMg8nxktabWnolg7E8G0sxmOLO5sqrx/OCnJ/zBCLT2Xqmf
1jl5TmVX11HZZYkuyvX1AQGMZhlxMQ0WViAyZSmLZ+4ZyT0/CTys0ML8PNNfLZby0t57SBKQtd7f
NAAYhLTWZ1Xow7A1ylmpkOZTPtBk1wOvzgmnjm//qiz/spZlvC9ofnky8zlCMcXGld2y3axzYzSE
Z0Fau49PVPtHKccDXwN9X2aOgITqXI2ztm+i/qTIx7nvUujXDQKoK9CFGG5mhW/sES6tt/B51wMP
PwmbM5s7gnGEOSUOJxP6SENunxZ/6hOybhaHVGnUoM0ODX3q5I7bignCFzllwy9C98h3iMw/UXnR
nXbAltK7gfHjaK2M7LCIbiMAStcm52jIpn7nHzVcoeyYzg7mEpaLkmpVkQcVlCTddsw8M+BHU71O
fu1CruX7KNnsLDGmKUWVTdjaS4MkW+XcDCCOsEMEXIaV4p66XqggoC/T3famflJ5cS5gOJdjrZca
e9cO17eOExfEVCVnKiRKxs7vsy54Vb9iBnOjl97diarMlprbXDWUqbMcNNqc914G/rEcYFRTJPNY
4FvQfi895zCaHsfYm9rXIaooq4Yz1Cfei+N5OGfYNaTcnkB+QYR+5S5aebaALzZBJiUqW2FQjUt3
VKpEzK5salDdyktin7rOpIcvhpA3iz8sFHhRNG2dHocXATbfkGoEreKaKysYvDEMdTa6LF41qTy0
DwpOcEE3cqJ5q3PzwM7cdnXyfbV2ZJCz+xuYGyOYI1b/0a2h0w+XR+3TjYoPDQM8MBtxOPMF7lp4
fcKkbuC8sp2ImCKrE877BAW8PxThabTyMQk8nRIhz6yc9c7g6dvAnqABA+/wSDI7FwT3FQukTXkd
e6q4HkhYjERProqcifE+TxZiHPBwaZtPqJsDZLrza/+yPl3GRoXF0NVrDFPSllpkPJs5RpymSxDR
+1XZ52E1/hk/HfbPZAXmVNRo5I+XIk1ZKuy3OIFp64VFH80VA/Md1VkFpkJV2tAxGsDVJ0Nryxfh
GF2kUAcNqGCzjbKsnsqBP3eCaV+yJSEk/UqtvqhL1QqtXViRrJZZaMrhwwfsBtG9O4n8WU1ilFEh
d1WoRnWR4+hRPrtuuetg1/q5PBTFOjd/QslxW84vv+ufBlUgK72H7a60nviA1knAc5PjC27+9uE4
jypbr+YqkGla9o14KbKKTaEbUNbrtgQJ7A4Ilf9UC0TJNLxv+IGma5aAjKC6LfoNyg4rfs8EWLR1
YnLyg54vXIRxoY/HJSuhqRxqsYIcU+5yYLH8EP9Q4FB4PbGgKLc84a3KTSycOM2nEmpjhW/Qm+N5
ECvK5f3JW+5ofI0NKXTH4AJooeCSSkvOgggk+1uSsi6HbKqg3MwUYzqy1PpNfUcQFtIoahd28gsB
fQyXTWyP5cmmgF7FkFfgX97PtL03suwTAFUfk8QiLgNFslEh3fzMPc7pfAT5/QZ16ow5C0m4Bcbb
tASmas59+gs+Mlymmt7HqMNTdVbTLkkOtEBhLyJNpocKOSzJZkpOpYSVZVTVzYMuDWaMaVSiDK+O
7KUnxoSHXi0AuIhXuJLcjPE6Hhz3dzzwVflMiYBSC3FzaM7qCma++EtW3gFQglVc2YS9yX+SeYa7
Em+kw47ek/aOzt41z43/frmJ5m2Hffqkndla8z1VS316+QPjWoAB8IMI8MzjUNlmVoybi0nPG9aI
45aq4tvxD0TX/nwzpZ226LgIaSFvZq6uAM8MxyToc8yHpLybhjG+8YCPXiQCGz0xn+bBlHlECoeX
6IFknx0ZCqEqv6EatJ/CBaXWsvGPeqatoMUWuThS5zdA0tty3rzOTDROe1dq6UPbl1RdlspF+0Oh
7HxyumErO1ubCORoXNqJ+iy+Xs1KxuOtXPssT141sGPePh2r/N8hE93wS90Std0Qx7xW4R/MTEs2
D2Ff9zFC9tRy1da30ch+5TBs4Qk03Ia3mbqxQwQuHkE4ts5GhquYMWzDbnRYM+d9PfOSHK1Vx90E
EHoktT6OsLKulEivQ5WXcOWAC2c6qmerCdVN3noLlHieZ6/vkDrTEG2GK2ReUrveoUjXhvC74Z0L
5+vjiCbO5PsN7YKWGbWPY5fi0lOsPdFN1QDw4/RI1owfpGDq9YPvKPLKO9c4Y+jdFsC50CDtSzTr
fBEGtXDFOwJfb9DNBkFhAq2n69tq/dvL4y7sHxcqmbNpRqqyn6OJtH73Aon1hOpb05qltKtkiEzm
bMB1WY+kO/U8yAZF+7LNpOffgJ8qRNCrzPmbq5r6DDIdPjjtdp75gpGEd0RrfITwI32tYyJSjBEW
7QjTWAcaDmSnrXyUOYiKTttXo2Fgf4vxXzMRsrjgVxeKyow4fAgK9okERZvMM1MBo2Pb5uyCkKqN
y7dc1lTl8+ZiiqKmn8mQyAE38fM11IPotknVNkp0Z5ATLyDDiayap9BmcjxXV5GPxvotq54Qb+52
Y3oz42wWWxdLrBvshTb6G0MtKiDOEIlTfkA47VtLJC/qY0f5uvsJabUXUD6ksGeHhQxMj01t6Z+q
Yy6iMl3yZQ0nm99/nyw8pLjdPMoY+JvGZLliiVmCOZFFHqsn+1zlJdkhI0tqYsgjy8+yRygkVIb+
NQVRHD+JCm+M5dPW1OXVfmHBbVgPxjYr48TNdaVfbdiPiEBNyl9MGz2wgofj23Aany2g8HdGgjQY
pUyTLWazMSrRzAmDV1BdFxzuVk79SCzge+CiVLGf+gmKQ2OM0xfejavnvMG1oIQl5B6/h1UjgjSi
4KD81IR2g/y/QS78cSSpi8WPGFXG9No8Ddcxse9x43F22jVk94S9lePRl+wOJ2Zlv2cnF3WRW6eL
Gm/hhZgN0ISf7mRn6Byt99+H++8ujTtK0ubKlFmepUaK6bOlIlfjnCBh0MfMS65wWRYj11KswwRU
wEMkNplpiCUSvWPvDA/5mnCQvXu6Q1s0lQCcCkPFTkGfkWVk3pvHjqxQ18LeQbohohjP+TvdDXkw
oAcBrFDyVog7EJKla3MHEiMbwut0tFLF66lnfiTyoJ9EqM1NRQBPGRm86+7Bw016kRdUPq3fFZih
jnoEN7NbwqPna3H9pJtlTR9ZPux8lDdbYhkwgK5mUhh58vJtULgdQe55abdQgp+f0meF7tKU93HO
VJCPwID1ZNRyChG55qCD82CP2vGUvCeBw/QcIbH+UYqDpvIXg9+Pa+v8phe2ZpHI3CCTm+R7BMFl
vW+vwTqxxnLi05dYhkIhNizqQN440mS8L6hIqV0Ep1l0J+JcmSsJAy9jfciCIeEXnOtnpSsffuqw
kyDToPP0is7/ZgdByrWPPw9aho9SH01rp4ssnQMyuy/32t2MgoktT0UHVKjcFl2t/kn3UMzPCgVT
2a1ynZIiI2P1g8mpUjjPb2KA0Jekhkbi0UMplE7LfRxjeHcR80ucpx9iMIzmHvV4YY3YopJd4gf/
GAVio7gcX5CrcLXZERpypwzLF//mW/VnbYjLnz3lPsCA2BZHaW3TLTJITZ/TsI+xILvNNEQLlXjl
09zp/JfRFLzlYU2OMoOEvR3YZpSnUWhXOaOPJTgM1G/Ao7qSm+FqepC1miXNqCZ1vwF05c86b127
s9TAZn5bavbontBhIR3rYKIwpAgVZLJzIrL5xDwRua375URDlZfaTxQQxSr76gE+H65iRfzq5r1/
V/qhXRnqWiBPggIQ5FLMqQdjE2W1UTbTbQitpvfLGdGxkaMH+f6Dff1kzPibIC55d+zWpVsCEoEj
N4ftw/4lFO5Rgg5k4N59C6gMLuh44jqjgKN6Y7TvZH0fD/w5e3lEHA2ezAjCGsHxCYtgPfZPoaCt
+Nwftoh7/6R09vEnlSxi19A927LtxUkcxn7kt0I32HaJhXmlhlsEeasYov4q9mMbqLpGgpw+o6Z1
it7SgWCFWVKYz6jIqkFSDIVMVdhCd4b7tbDRYDJ1nJ0etFvpykcDv6FEvpv0lPkWuAMeJ8EA1V46
G0tGN2WXakrXFRG5qM8SN0yeplz49dhKJ/DH0GI2VzhsLI6gh6m1WZ9FJ2lXNlPPctcHiGGTc2th
1DeSxH9Wku0mtDvwPh19Tj7dwu1aoUGYAXaZTv5RG528ANEzAWi5CrJ/Fg6to4jdqu5P1iVpgjvd
wUufgnEMFlReSJ7gIxFAjDT+Kj/1Eh4S4mXg6vE7DtPzarzEryWiOv/+VL6wTGXFoExakf1WJ1c5
c+pM01icmVdEd71G1RFbZv1HxOst+vkkupy8yV1mGpzd7tjr1DVjYRii5nQGTfWGb0czVZBuZgu6
DABiBfKVR7fHPW3toGWNO1IB4keYCBi9gwjI0m7nYinmfbvFIqgat2pMVWqV6pliaJRQjbJfHVUT
FoZlCC2aWztQ8/Ef8k+73Y452GJ7up6WkFwshLQYbmGXGziBskhU4LqqSc+5u53KLsqqJCqb+iyw
CBYBALZ6XvpiYpJnCwnWMR5dEbZP34ebzGwYKNEXDQtz3moAHBL9lsZaW8wUMOuqzGBL/bTh/Sl2
ti0rTf4uum3Hu4oEcFIIb6we0lUsLtTjZJ4iUvSxRgBFi1JAnCKI+xvANz2pGoeFXEdf+30/z4/C
JicMJ2/so4Ooh/rB5k2zB0J7mE5yrBFS1MWXUD6gf4rly7kShYpeo4wlAJNSfbvROhCFNW5ejRFa
DsTpfFIvFwE8j0O4belJ6or1QZm9fmUcibKSISYkDrwf6YosM0dVO8WNIyAt5NjCbUal1gJvdtQT
LFgr6XAn5jei16Npz5P0LGrjDHI25vjFXQE0dLfFZ07IYIBH+YmUSG074vykijokT0IV8wWd4jZH
k92sk0iLWvJMQ3lkm5WmSlJ2bTlS8Djq9D0LpDa2ovV8tAsP69H4ms9eVBubd3PshogRyRnJMtzp
QELQT332QM7uKobYzjaZxUD8I8ly5QgIgf8BNFgvMaQrjAKO0+19DSUt6UNx4oly3RyrnM/GXWkk
HeslIbTf0NV0LPe0rL7kvllh9ymeS1a5UfTjWquU4u80Tf53HTIq8GmOO+LyxmGpeXfEqgK9aY8L
p17AahDPxdAnNNGffFdDx1w1EZXEliIoTy2eMHppoz8WJf9hn9mG0K9SxwW/WF0IBEaguWq0RLzg
ryHbtD+l38Pb/JsnqEklp7jRwBgCMlVSP1qpPBEFZJv+iXZTL9lmKk8qKA0DE0BKq0PcSDqeS/gJ
MKomlzSs7l7FqhvQD/BQbCX3S4ThzIjpiTmIOg5VpxbYOutKS7Q7ZinGtsg/ldu+/WaS7R/M0bvo
/BaB0AL7RmBcIjl761LpT5B1EchWaosoH4ejlVaFy1bmCOoJ19lPkn9g7BZ6jUZXisgM4yqTr9mT
s6Ypb9mELhDjqMo8RPjf0M7eIbZ9edEOycucwYMdHaiF87u7RIYjapSLMtny+szQer9SKcLM/VUK
Ge8IlJfS2ycsR+6JkL59+1Sb0SpoqYrN54LwB3KSD5c8ucVXcwbzlZBx07WyhSkr8Ewl98LpjFwq
gO4twYI7Hs+AuvCTanbnvd+sJMGG2jv3QS9gH6KAArbdHOSVjN1QKwD3fI50p9J8/6j8/dvJxycp
DGImaHV1tDlqKTaH9LgHXrNYGzPgLiFQYHie0+eF2LjOYu7HZXF1suoEuXN20Y2WLJ56e7ngM+S6
IaYPMvI1bkvWc2BXwkZEgo4mVZvCuhr/S1S3XG0j65uzvRppdwoSoEiy5JPZ5UVHohWH1g2qstV9
S3/mGC2EFfnEIpHpld+PRKqzS86RR82J5HDug5zODJ4jt56U6QR446ZEtCVqNkLdKzJhyO/sc3n9
aNcSP80FGtJvA1VbSrDIGJX7v6bBqUZRsA+qnp+0Nfq8PexOMupjysbmZLBuRIw7yv2/+3GWhui6
+6dJ+dvKCHg/xW68OXJKV0j8lq3kN7lSpsxm+0z9Ai7Omt5scolvgkZ2qRKn1uhWLx1sxS/N4HZz
uGX/81PWTZz9d/Ki30NH5vSo9hH1yohXPowq0Rqd1HDA3poMkxfDynzopBx7vBGFHQX6nL6suclQ
vhoU0cISbgNdCvXcQU496U1lr/8xoJitM2oUkZAapErC1aOuMjbo5Ni7Izm1ZUwmfAQXCoJcfPeq
hqI/fzUuKWulEPEvpdxSnbweffFxN15KQozYlZaLz4liMeWwX2RtHrsEGqHw4v6j6BUwXu7SE7KC
PeonWmlONyZSMTKlp+n5sWd6ef2mYt87eG8bJiPvsy1Q2NnwgjgePLIi6pahl9QQUltjdoyIPSHV
r1h5rXJNUJKBnMqaUa13H1v+eHo13pC78nn9G8/rQsw6Hjimm/dnDOqWdjAGlXwyrNC9qiVHLK5E
L2lKCBK66D6u7o93d4rKdMVFwshivJkN9/+t9hCDkzUwqi9GmGj5jRa9uo4w+YLokfoWNQIbWR8M
HL9ki/SkMZOCmX1Z23dJI6/z+U+uGAe3UH5toY524KNSK177jp3KTmeFhD9+iQDbJ8BpMc49uMPv
UUSNEihC4MxVjb8iY4XDhxMLgNiG4VjSjZZEx2I2ENuJrFzhaKQ2QSzxkgZbP78emcwbfkrP4tUh
T+zzMTVbWdiol/PG14eVKWbhQ2rSArNiNeUUE3f9GFxP3Kcw5Vqcu6FsntcUZQi9NCJc7yJkiYf3
+ohtZVuRnAsVKkqkzlJUjDmYba7KWv5cvAXudoKa0EndPTxx9dJEoROUmGdg+p3HIzOKXPV0ZaYe
6S/Ve8wcJnNAJv0EqUWIiIG7VT0l8oxVUC3BxxVc+qSCGz0qIKXPAVLHIh/3GnjTeuZBxcINHU6g
NuEkqYKUq/MxJre6oKe6mQvtjHKsrKbCsRKrkroIEBqz5TyihrcKk1QehvY8v/zVJXl8+OsGo+z6
7K5OfdPKNZflCd0AM51+RxvEjuFuOQKIVBipWCBJF0AWVeQKx4mJfYIP/q0qx/aYRGrziT65YbFZ
iWEm7jxfm8/oeLN10qXWunisWvq4v9YjDum6/dVEdmmZcZS5Fc2K0vXaunFonU/p5cdkGh9AgkpX
5pO6XfhjXEoqP1E+AtC+pZr1WF9qcxD7ju55I9huke/gGefLnKg94sebm2kQscYrmVY6K+auv7Nc
XQXgtn4cv+U/p1QuazQLWgIB4eh8p/YCncZZmyiaYRMFKVK8/xXmt0FM3eHjOoiC8u7ItHVuwbUd
FVEILow7X0Khh2P4F9gab/cuBW6tKEEXP947dsdt5soPGMnVUWTn5fuNvoc02h3Wc48904xWBRif
JWiiL9KtnLVrJH1rFczf6EUlMDS1BNURry8NWUi2uqZhWSyNkJUwXLY77eaFbyxU4dj+ynsP2ycB
4d1zUmed4WpR7QSvmeEwKeaUYCdRGmmpV0Argx+FaTjQBd44HIMM4WJt+qbzXGEf5Vfb3+5o/mHV
tuHSmfE0Fgz5knmiHjkm+ZFLkDa+AfhWy0LJQN+0DuGuNsGy0TYAqJsVfB+pUrHEEA5ddCn3iy0v
uapSY1LHjyA4iDaj3pbpdvEIQg5uVNoKrJKoaBU4PRgbvc974j7vlD3ykSHhpioTRHIeAgeFEeDQ
/85bOv8gsHrr8C7GSX0Zc16PuknqCDdOIdopcKBKduWHymyI4f2juyLCWAyGSUghhQuEPO7WcdEj
2s0cjabrMMPQBcu4Mxme5UCPmTJsSGIKGHm6us+4SOs87ow5JNgEh57umA4W3Ec93Vml503937a1
sp0zxEXxGHT7714+DP0uS8jRuFSVhIRDwcFYjeXkxBMG9PnCQnYllgf6oC+QIQ4osnUWR38Av9Kp
QmNrkUDs3bXF20u8En+jGK16zJPZ+wt8PTOJFMPe4XDuoCKu3WUvpwz8acu33t3JfLN99L2xMgdp
HW53xuhHXC4QAMesjOdh6UdHyeUDFw/Z4pYx6COWYso8nP4h5yIg+pMf3PWxaN4uETGZ7Dn52Pa1
vmrX9+Mx+0hjjFUK3Ui450D1GeaVOvM9GFiAPgI2sioIvX3ibggvnZef1osrsaL757v3eZaSaWuL
H9/RXkh8rSzcT/OeE7Tx6UmQ3dTCLsgQOO9KusBSrtRE/P9Itt8Bz0jQ/IR0pbv1Ua8bm9KlRF1Q
irWMW/hezSz1ta+uNa9n3vaSwWucEaHSoN7ECMQ0ER1O+YNlFyFaNrSpz6EgRRutoGYo860XG90b
A/rSqNHoqPXO6sC/7kyQBStkFp/8SLPYm0T2mkxyz1UPfT8knI4EZedOqUORNacwsf/1HYQ9aX5v
aukcGAFE5+rHBE/Mx1zQyz7bFSqZmLKmLSA1CudJOioGvSNuIJMrm1i539+WObvIpTYod+v4YN6l
UTkDpWN8f+pvErrLU5TtDEh7sj+4efFT/OYdC2rJYi74XzzeIz71ZpIw4aVJ2DwT/vTY+uPHqi0T
U92V7rcWF6iWUtPTIKsIA3ml2N/zp/LRx2xxkefhIki9AXShrGiiIgTC2GDZwHBHNap1Pb8dfpT/
gO6rsYp9LWUySf52p9zu/Eq1o3dMHkKuz3qqndpr4iHEEuTvTz5eRPFYlsnRGRM6RL8ChvYckCl5
YxmhvD1Xyf7KynRXhMIYh2fPOm75lwBVAsqHHCZDnaZtxL+vzAOuLwRnuoHXMwvj8HUXmt2TkmgV
y4DjjV6nQkySd9Ozbsfx+snKUKRMiAK8GZQJHxaudhzvE4Fcs0WaHuA5Sdu8li2PW3qMGzratigv
ZufX58gmQmKc20WP/EdfGsAmMgk2UthY/Sh72GbVOUHulUp/oCL7gNHN0D6w56jP5jNetMNZfKj+
8yOwPoazZaiT/yuwasCf1FUeC9IeRbpxhn6PZuQ2KCtH/3rkimNDJCXUt70pJGAb9pWCKDU26qsL
A3M7Kq67TI1GhOhaHuie4sAIHq8aLLdhEN9vnchKCUosPGQdQI3PIx1USb1Oj40e9D2JWfCObmU/
5302GWKfn1Cwq63hphReAVmbDEGFzLmHCXlhpQITCo+eoIDsN9NYoAnryeITVUfCk/fuwMOfCyax
GNVrpXkg7bhuhoMwEtwz1Wiz5j2xwH4A/goRY+4tG0rMupkrXdyQ4Afpmsxh/e/awknFCTuQKCQ2
x4XZ8uhBgddZh2oJfYNW+4oIIhnj2v+eRkZmBD/a99IPHNI/q5uxO0LAfW0VP4TCbvzSIX2cxylr
xNpF9SDfxzni2cf/DNOPKTTPIKhX2F3hbJ4uuE9paIO9UxASnGr7m2C9cnc08xoy3IB3vsqHrL7/
syb8cdsWxYip7A4waKW4MLJeifDc7j2Y40/yQ+W8qqKNPQ220+R6dank1sr/QLZtrpEh/yCAJWph
XF2yHpFGumt3vNLRRK8/J+J0Nd311oHTFlu92hC3mUURLgvIPqGc9E0Hqj1iHxjDrv8YVAly+WxF
L9I+iBixAR1kDKawwXvihtt4iRNtDOMQ+/dg7+Jwj4OZDiRiMu8sGxSDKLf4FX+Hp+T9xVCWzE4c
rXGzkXk9bRwwxiNqHbK9E3MkqLmlTmHDSWhn1+4UMjjrAPJz9JEAeC/gA/logXOeDzQoCibc2Pz1
YFKJdukBHFhWY1GBOB/5NgzmyJWbAffEzYFVroQFavMXzwYdmJogsk27YxzBlIGiWvZgHHBB64ON
Q1YcFGoOUcwmDlUJtkZ/Qkvzxg4YRhw03f/CDTgwOF64BlolBCR5gnyA37mQ1qSwoK8inx30Umu1
Pc3LgW5cXy3eIPzFGaohh2SOI9agaEVu0e91xXQmDHHf96L97kDccxXKr2A//PtJx/5euITDazvi
wqdgwn9gymg04OCbYJhQIZqmHlYLffawVtCvgso9RLitNNbs8COSF5DimltdJHLoVa8t8f1YGUVg
hbhrWXYPQMZDlSFHonzYRGjwgVl5aPufaCvuajV5i7txvAU5ntK5B46bdiA9Cd4XIw6YUf1Rk2+q
6exIPpDNgqr61xweJ6ZIt9H6i3DS6tqaRXTgZZiXj7DyvqPxep8OKrHD5eeBm2T4NNHoJP7DBj/y
WGPHwAAB1Wtf6FNybsEX3aDfIV3Jp+tLTkh7/dispWVx/Fto/8JhfTB7yWXi5Hybpsg+mguUu9nI
TkDNeNdQRHYSIcAyocPmDu3Nj4YoP14D++u0Dh6oOUWUdb6+Ab62JdfFnlPkAwXsi20KKuiCS+ut
0ijO9HELeiuhrMUDSCf2qSG5BjT3Rp/fNCbKZp1OyYajVVudhzmN7NJ3G3wjWI9eyPsxMdl35f2G
JETFrq+SBBkYMI+YCeL15obfgedcAh23A+nUdXw9D1ClWJq0CaK7pg8pwW73Im7E2B083Xd71LLQ
8c6/z915/mhQvmtO2JCkOtWBDuw4EUWC3KZnm/eflp4v9DV8ymfcrOu1BrSX9XxX5UchK5j6xOGa
/TYsOabH1NLGsMcVozUxvUZ1hhgxALektUvTjBqVXHMO77TvC6EjQsmSkesDWX5Q1cgpRxK21gK3
QnmX+wmTNgl97n1MEiUMN7pXlha440dqXYHAX+ehfij0wQPzVXzSqzaj/d+TQbjCCmeMLlbAGlkr
HJyflDW4whAUrUjQapejdAor8cttGt1YxcOzL11hPsdBTu0KDNjILURUoCjN0s+KbN+cRjVmQRGQ
VJfS5reyDiBJ5VVsxMJpsGD6wnriLaZGmvTBnbnDpgwh+ib9FbM7n25i9vc1qfrcjeU4VHO7b9SG
ERzurcqKAZhdnGHQaSMPgmBQsmX99U9bVQlXt5GlKFqADEeVTIZAULWWdhxrEXDl84mGNhP6QRCN
kBugEca8wBVBLhK2UqPz7UViWhSLM7GgBqfyyhGG7yeI2rtHbiDWqpfV2NaIhR5HMMZqeV/+XkUf
Ya17WzQtFfbgPpfF1qX6AkbUOzrRtCrABEC63GHRe6GEPQq660UTc/rtU3q+YBbJ8vEHW9tD2cFi
deVAAM5mVktsM8s4wIzlzOytBvKzOrldOyvJt1PYOMsfoON2Rzcm8vyfOH1LlPdpAJ3fr8yUXGNh
Fhem0LBppPpfNLn/VQwDvGv9rXOjNkR4J1ob0HNwplFgdnDctcuHlk51O2qk3aTVFruYNG0m6Nh/
ETq4hwogEmhQKaG9E7iu64WN2d+Mtu/bnPtlNp9x3Ad/TL6SxInnGQbvuKv6I0x8VDrWrHUiY20x
wY+Y0oEaMR2sO01/6l8S1Nd69iS/dDshFvGx9giOTZFTcGCQSY3J6IFG5ZRnux9p4V3FwoiqRiye
x9hBvk03bKVlKRLZOCLIWjSNVuucuU4e9qobX2URrJU6XqLyBTF3AzOYm+KDniApHRj09ObUgthO
K53bzI2V9OBz3nvVu+9Xrjlg2xtQm5QsJQaeGcrCmLVmDnLotQdgxYJEzDitqDqrEcmAD26JVxIl
3889wW5Q820S9Kf9yU/JZ986Q0608rKZuVJq0kVLx8jol3zi79MzGwG485VWE1hzSeugV0iLO99D
gGHjXlX+l4aTcZGPO6wXXrhEfiWG5+d3VKsm9y9qVeQt4EXM/0aIL47KB1Nhw0923VAsqLAySd7w
xmZl9PRhWfo9Hz8s/1nQ02LV0smDtKEj9NeoztA2nAVwfJTVy7ScHxMwNcMCOqtSut/UrXtfykBs
qTUW79rLK1JSCX9fklaSNayc/P1OTZHaOqdK3JRyB8WsSYXaYI+zSlJOCxSRRZ6oM+uGKBMwU2WC
PCzl4qFVCSZaUG+7w6N/v1Q5dK98fr9jKHpZjoUzI5HuCNnEiRBDTJtgKdyNODnOrwgRZ4rgiT1i
QwGYaQQfwLCdp9X+J2u0pN8eUVltFQYGTgdm0tdhckGVCmWZyBDNl4F7kKINA0fOEnToF1qUhA3p
+0YpygPwLok1M75LU9OFG+5NfLA18F6s2yyRHENyZAP8I3TDVL/gJtZc9r3vIl/u/H9aHWCETOfx
X/2tuZzWKoWebN1vVEhrvlNnm95oJUSFsGg4fTFl2+exihXJO2h/FsxbtPhs6Ns2KnTrEC36STig
mykA7/AB39ceCYD0kL8zZEPCjTaE/xTiNGgKHRRl9RQ1Rdpoi3HIPXSR7VIsUFRH+k0KGr6+xENZ
8eYjgqdEF94VQHbmC0TeSrHUAomXUmjbF8jbTPrbqN6pdbFnd3R2P2CMCXJLLwmZeNqrnbRC/5V5
63BmjtohATiqB3Cja3aiTj4z6fK22zqn92FuuD04ly3ixP0A+f0yXgtED7U7UUz0/Sz0dYR/S2YT
CzgIrZNfiqqpmOySQ+T5FbLAUfl+RDQ83itgd22cUUFcK4iaLVuXQZNZU0i09+eEPZKj10QcVnvV
v9e3o9Yz1K3X745Uwt9+mA/SQmKqdaDTR3SFBgMZ8Yu3Udje5TY346VwxF197cQUFmFYcKN2UxR9
5LcdbVsB6MGySRiX9+6cGHez+4G1Qd25qwop1CF8HddpiTDp0GIjr4Uzh9jstXFSvpIek2YQy8p4
i2TQPeQIMLB9n+JP5tOkq6MnBrd1qD3nBJegWVdX4LrPUceHfcPN8enSLZfxCM3Sa2bRYaGquW7n
T/U4tpMCsK3x9kk5HWll/ipjg9Y00NEO6R3uVWbrnsKIRhoiaKF+L/TTWdcaOSeXpGxi9YdHhr8/
xH2wls1d8B6N0ECLFMJUBq8mplPN9ZsCFEf1vrj0dBB5Nomu4TYCYesA/tnLWH08TczQJHXXrZ+z
XIC6diLLeAMavVzNqyHuSgmDBH4Pt1sfHW+YJAFe5hD8oqHsEmJIQ2VCn+cg7v+x5O1AInERIHW7
jcZXADS7VkhkWjTlpkzjyadO21NvJ3S6IcO37VmCdaMLbaZ+6UHvx7oaZO8I5OXxAd5ATAvstEbS
qTTxVIca2UuN1fzZFA7XI46DM0wroPWZRauY/Ce15WCZxorO1j9bmqv6h9zYrPRZp29HhYhiiaE7
bn+Br59YsdFPEpcrt9XOG+uyndCeKx8ufXlVUVnNdw+ZUl5DLyvjDog7Z2ZXwDYiPuRzsCjjpPLL
3wo42dVfVdlwP+HHELmghapUzava5SgNRi8ry27n7UTuLcZGmMEIrK/4s8AVEE4rf0ZMe46lUtJi
jq4YZgV5ZG0W12L3MloetIr7I2XrjCXeULpnee8uWmKDeTeFYVAj/YJmVXmlWZ5Wc/8QzmLlUj3i
jdsRYgCESUua7OXRlbzS0kG7CDLSY/+W75TKhM0gRkl2uFDuWJk9mitX3eZE9OL0jHkNc9koQtT6
BPAHgxbbMGr1ZeaM5e0L2nQ+G17FAS7OeGq5wIINAh1a0cZF7vPCKt5Sx7I5Zq4smNpgz8Y3G9sg
cVuBtgmdP3onYntBcBYRn58c3iUB/93nPjNke5VKcQN4hYzAcwcibB8VP0Ykksz1rBCwCGgLD5aJ
ullsc4L+c16J8oJb6bgPF5WF54X3wlo0w+yz3UAYhp0mLxEm/fCXLkKnRy4d0yp4QZH5KgycS6NQ
VKf5DiMKxGj6VNq55Q32fuWy8cEMVVmlVdQ6j/nUzuzcWGFv+pUkELKLlOmryqp64+3VsQZkylED
Q1O6KJDeRqVVNn7cAegtx9HyfjLdNLhqa7upNGcIdAVQRmfA1WVOn8jsSqchrNkk8B2BdTjuHNlE
PQSJaYw2d59ZIhibU5JPaLmMhsLpW9kCXPjeZGe2MKrceigiHARkFdikC3Tvh4mdoGFsaD5MKVHW
tTahB4LQfIbxil6SrkT0YlWu6zP5o36taG+leATNqh89ZZS7MElR184Jvz9J2q7XEujATBEV4L3C
vAmVq9UEyg84s/i6ZeUvo/A+Z3x9NC+f0DL76TehcjvBo0jBwMs/Rk64AfCpz5Y7i6CIqRcjRdpb
naFRYDeIS2wThINj0h1j/7VwfqSagQkcPZ7zaURMRuwZuR3LRIQZwrLUm8nXpElKdsQuUC40ZKU/
8OLfOHo0WeJu+MwKL9Cx3gQgre1Ss2lXXy2P03L8/fRhrAxEiSPEdOe5DQ1L74/wumGxckvzXltG
y3NHv4GAH0cQFWZJQiYwarWbuk980nq4Cy8FRIMnZ79tIGfZemjxxuRzxVG5eZ3StGfPBQz6KWv1
UtIBxTBMTghKC6Q1aqXlxHNz3xCKKGa+vpKUN2mRvGCKfsV3oxrxeVxYuIG6Zoe8dG3a8i40lvO9
NZ3C4BXCDBZVYkyVy+ESlXVh6r7n8+4jRhpIDAqf35OSZ5B8oOqdEWg+iwk0KRMAZLA/p2+sgaZa
ifawEvpI3yAdg5G4Vfen723rZKLnfblExvo9GQxlInAjsOWutZp0peX3Uf2eSLDc5upPJy/uIWtY
n3c3WzyzFHpP2jARuSW/lnZ1XvBZG4NWNqa7Cj5tb0CIPzen8myItQD5yajwBhIG6zHxFhNdDFu2
6v5jp34sNgH/jQ+oD0OvYEIJG32VmCz/Bc0X6CNV4PdHOfEguV65ZrfMVdW38A49xli2FpkZp1h4
a9kYsNpO4x8vbgsPYGYL/jCKOYitedbqS63cFsFg9riXtdMFRkPdpESiab6F5NXlbLRMjnOMs1WG
oQkG/P2gDTu1jEyOPmUoJl7x84D2c7YNGNVeT+rzAdYxdpT+/npTFSa+nn/+hrTefglgcRfynPsm
P0V3W5evo1TStFIbX1nW8e7QEUCnnu5u4hAbI7VgYMt0J3yB1bDibdl09p4y0EJzwsbN6hl1wRB4
+KPrMO33QSMnhIIjkgIFy5x24vYA18ITQ0tVkLZM9J4SFKxmfwlteSJlrR21YGstjZPyjhcVCKg5
Cg6aRxULT2QNkV6e4g586OucvaUQWw1du2VddSvUdgbDuAQze/apBR6rdo+RIQiqFAfrX752aGKZ
GkoMHd2WWfHVnBsBaY+9p1ANbFucaHT6/cOKfUuZuj8v9jvasdlVeeZmw0EhKwtCqrsyTxyDcV/j
awNVIPSVzUsuONFustu/UCRfR7p4yOtMnWfana4rcdoem5rCRfUR+c/wxOhE8rpIELVDgUi4JD+/
Q/IZvRNHw9NCJQFPnbWRxe34pezQlVb1EYUq40//cvM55KEI1ZhZep08KZ1l3MuOCqWFPVajKxWf
E5e9k3IFhxFzYaKy/WDT/uTh3MGh5QSXNAaXXa5LjZQTGUXZHoB+DsIigwU43urLM+kAW9NAQSrT
GgQ3N2lylp8YzEc25lAuxAlrvYgYfI2L7i5pb1yaFcxGgvBR6od9bJ59Dblge/I7rxGivfepahNm
56tBlUF35H7nYw9MTO+HtBf8SMGUpjVb9/vMkS9h41K1xsVaNmzgq+iywVjg5di4zK/U4H7FgSRE
RPX/EmOa81gDCc/kSDTox/FMHHGTVOPJd4ezJLbaZZ67wvmjeOr0z1Op7Ycj+8MRdIUA1v0hHwzW
lkuRWxWBvAK8tQn3a23jaip46vyMIgmsndE0lV3l0lIthspFz3Fayx9uXWAtubGqv8afMp+QW7ZW
db2nesiEz9bO/ITPSl8C4ok1defk4c7UjgeD3UucgfPD2bWCcskr93eqHPyswfrie/M6HOWoL2hS
zrJV8WVHwqylD23kOpcnrpI3weJLcmF5wlEJN1IiRmYj2kQTvEyC+Bi+rdMUJoPpwbU2WQcPNA6l
5FzUnLrFskVUy5hG0jI6W3FWXtrD6DwPBcpPe68zUl6TfnCBNkrauoh3TMP+q9m/h7S+tHUDQNw/
2Y/3C5+3sJd/wZHvW+Cy6uciiL35SEcnbGA2FgDj3FBvIWYpp4IT51S+m/PHwV7wWlQ0vQlQObQY
bEesQ/0Mtir8vBfm7FIoHS/iBZ1UY5pSJCm8UwN2phbKLU/zLmcMLoZ9vUiWtQn7YKGUW3Fue+sx
mwk27IA81BPlD1lptla2Q2Z8g1RlAv4BV8HV8lfdPIiPwc0XEX3Q+l9B2KUC7dyzYblXqJojzXf5
u2AvrKO8YyVkieLEKicz3lKubR3j6X+HEM7CTN5xChC1068n/hXHAbqgdtdvOQYVsgmjDaz1oTCm
W0Xx+9qPdsGXURAa18e+YKhlPbyO23n2YZlA2uKJRWi1s8x6/jlHzioh7blK4hkJxNfPEfQVnb2Y
9jK5uxXEWMxNFUbrVBZiaW6XrHcRmDdlrCAGb2pbYGBji/hEKoTgDixRCuWrpKs0r2dTWLgH1vik
JaQqtGMeLLQIYc0Mm60/aSQqm1hgT8QqEjbi5pbk0Sh0u4rdDeJtfdfNQjpCkP2gCYMvlyOsOtZ/
k+tllkYpsr6Mz2PT4+fmP7v15kUX6aufRtCTz1oLSjg/rMob5TaRYCHZT8lmmF9dJqepV8mQ5JZE
q5rPDzr4MjHFzezuEDPTlO14z6ss4gGJzBUovGyqBZX74kdTdsypT1+BmxPF1BAsJjsORXanrjXv
Q2QZ6ottHKAS3vABJQO5iTscWKg/T2XFa5RJxWtsw29T9ipXNbomCiY4oQOa9KyCLzBUkOGYB94e
odjNdZtEi2ldRTMJtTAkwFHeiM5IrjN9iQ4AvyK8UPnv8IkKZ//4ChG7pBDjgudYhK5QhL5jkglQ
f3B1X5uZ7o4HQ2FijGBQm/jOzn0bx6czci9BqEu26Gc3txqieip1v2S+/FOvZWQukN7/YZZ14zv/
QOWSKAu68Bx7PhuvmTqXdn+P357CnsvdA4D+66s/IaAFM14Qn0efl+PIQldyiMSdYd8DBMX7Ktp0
VxDjM6PUvL+qaMQJQMQldTr+Njy2Op2mSjzJcqc5l0nzbDN5rgDQYbQtmQ5LLAy5enifz+4k06r5
y+sYH1K+0WqntzYi7vdPTSP1+Dy0O2bwmyNxbDEFD2Wa+2gddULmQAO2Xj2qsni2zLSVApw5jwDw
CBpsQieaGPDO9eEZ5VjlpOqVSLC/m+FBC87JbPoyXAqqK+SafyFMpEqKi+aMOZhEzH3guTTXm/cy
vxUGjgC4XAyoe5IVclBHYp4S6jHz7x7czMs1lVycyEIYqpxKEnIQaI+BxLo/IYZeHE37ZTiFkq+X
fqC71eM+y/5y3qAcji+REHs8vuV4l3YInUooJof9E4QCWY8A6WfnY12Whgf1tQuC+jHYQ+RmolIX
YUzd85nk8uEyEwoALmAWXUfaZj3I73LhLbUuaOx8Hicwt8eHZicNsSWZTNMWcjCveA+ALcC4JhFx
961BVOZLfPFuirQXnQ35CgGKAKqBOgT13seDSXNtWQEIWcLlPsXHHBy2oYV1GWoOPp+pt44D038t
8Ncv3ltBkvAzhxHNdraGPKc5a32MJdNvBB2D/UQ35gGqCBSI5deA78HFJoOsrM/Y9Vzmc31rLUnT
IuFYdylHUzFviS7BWDHHrZtVgSGZ3hjRAoYItNzrOV9MFVROUlfC7xXBa3a8H0JqoGbyNSkLFGqq
VliVpLMHylAIT1jBb74BK5YPNXiAwsss+IYsqibwwMSPf8/U5fhTC/X2pFF0ZRr7m7msRcyGRT49
ff+BcHlzlP2GGUC7cv4yPcjacIDJLnCMS9uJrmaAIasSkMgUXg9PNyFNJMjXiR+Fd9D+WLt4E7/R
4XygiMNyod4otRmy/APT4vxpDq9Me8P7xnTLmv9H2TqG2fzpJq2cUCUIgELAxtyIm8sguCkiDPB4
je4jss/G/55xEy09dB2NT3IYU+Qn76LV0cTJdVlc0+Nv+c1E2WxK1IT+qKWPjlP/WTr4xcniOKRS
sDuqtrK9dxfvYkol9hb/ASCXwCSO3stVw+tMo0Tzo+PzCSaulKZTOuAF/RX0yWJo3Kc8gQn8PVBI
ljLF+I90bQ6mGGhOvLGwA1CBykGRzY6jaB7tSq7oX4YWnhhPbQ34s/awYTbIw2vkuzqN6uKPo8MZ
KL4pQgermnkOpp1DN+Aa9WGHW+Jq3kbjj6fCmGrtFiJ5y/xX4h9WQHLGu+6e4EfuUoMTdOMg5FWe
mXLQHtoByrL7UOuC/5sQ407i+PqAxrKH0Lk2zCSNsmg6twv2/C/sTsErCkGqUGWJwPtiFxMVoCt9
O2UW2ELq/Xab8tDRPUpd1ZSmHEBjmsJOMAnJqO5sa9mCXsL7lu1OE6a7Af00lKY1/E460nJPAq5r
s5NDYEVkIRZjfkkAe6aTvMxSzZtr6Mw7tASVOMrHwo6Shw+PjNsfo4fgocGMJIEY3uXUr79F9V/+
x8Bb7rBV4hy7f4Nq6LJ7lTbD8PtR4MgJSgaDATTQrJk5i45S8ioCZnVmtsPZhW20O1NSCgkt+/Sl
566856RWl0rlhxS+RldJvZp8fEOtpYxa+CxwBrlvxbu+3+iQY8F6tFDUVQ6aIbAqWOsxgYABrgnf
QMxuODPwwlb7D7vLJ2qrumy+wX/Y1y1jI+XIV05atskrYNhGiz6QbXeaGL9RNOa72I+mTt6UjKJ2
d8DayTr04qnzdZQLa4lVBk+mV5LJncQAqzuvU/ciBKlRnRdCrGS+2TdtstpbD14bB7bR+L4KnP8c
wBHx16zRE9Q7IJUYiAB5jZFraeYCxWJ5+gnEM3fShZZMpnCgEt2jt+gGIrei4bX0IWfiUWx7+M5Q
ZYH2hbCaFzfotC0SBrwOXFoCN8NhwCh3KYN1mcC28YLXdiag20Kdy0XwzyAgJVgVPn8oOwm+EYa/
VqkVazjnONum2aiG+G9pkBXe5gbk6o0pl8FiDnvW09ZLvM+cSejz7IzhK3ZWhzKEO9Qy7ll5q5ZG
pz8rzlV5KuZZgjNJAzXcI2j4rV1rQj2gcuCJ/nWrCeJNKJVfY1/FhO36jtHeojz0O513T9RaZp8/
9dlqLx2mOapMP2HlW1vpsWxlE6v9gRDWtyuA9//wEP6q5SByYC3SOLBT6C2Z3c8/qrL/2qNMJiGx
dwBrDLb3BwwLebNSJZZTo7M0C4yzgpKm5MCwi22XXnSuWEZKLFbduv9jgQDpTnZqesA6PeV6BZOG
DHGuNsSwrMChq68ePVnOvS3Zjd1ryH9TdHkx201guRvMZE8umwx7JzFWxr0ZTanpFn6C0EccA3n7
OmblrtoOX3quPeJMPotB4jIUNm09XWKGYgN6ZFOXS1XtZNevq+UbXCwyMEPm2EGcP72NyJ93YCHq
93qxY+PiZuoYHaW2MdaMoyd0dRx6CwBQBmwggml/OWqApCYLEfXG40yneOCMQ9oaTgnqz188Zn5O
iYyNHJnFwzRdSvsPi4cnmHJgb9Q84+zrdA4cS79fmj/vgYOfiCOLArCs0EOrcrK3I2cBNx82azwy
jUjj0Gila0eBf/jILhAHtmZO69GeMh0/MpQYTJDJuTeg+Q+7yQ84LcFxgnJB7gHkPgwCMg5jt0kq
WKbuMo2IdNoTGFZ7ns2dWcLg4VPSqJZGve8lAw+cYRrRcuYCBwcN1WOECckhcCi2ev2KWNcetWyA
tGu+/SoIqSLpgK2EBBErillJLvGLWss/vgrQ+U2QuaokSlMxQBzWGoafUJYYIDPmXaoS/O7BKJFF
8PEtKhYw30Kxh5R6mpGYPHKz5atOAQh3db4CRajuwtQICpybjTkgjIuXFxC+hoXoCESO7gJgMdEs
wHHR95r/rtGqsScZxRM48q/o/2BCwlmE2ESGSd1tzDwcc31lQo96WGTHk9fRGz/igAhtb4HrvFA0
jeASmEMthcQshPMdml7HpCkH2jmIQSCjvrcVRJ466hj7yzVkfz22zNit//l3EbRUVWTGmKAV5bXJ
bjfn74Wyuv5FxYklUUajM6Buq5aUc/es5pI5whPAdvZlA0Wyjhj9Olx1r9j/IYWKl9YLSlda60BN
nYnmyuchdMOHpf09l4YXKF9i2bMwJFITNZ4rfxw2Se3AJA9BTJe7KMJSfF4zznog58YcQIwCJ1aD
6OYelI0A17VDoffOyNcs97GNPMm8SA/ppe4Yhi5uxZo821iR4YI8AXj0ZkfUpH/QFZpyOCbP7L3T
E02EW/qfFY3Jr9CmTIh4MI6kSkYWyeRuk80VcziV5cv7+QmrdECdwH5bj3aluctJgnfRe6bF5P4E
CDUuDHZxAcr4ExIXdFlM7kA6LIe2DacqihjktSkpWmuOebsvsGUeH0+sZZCYXZRM+vBh91i2ibpU
MnPZdbbKpIQ94VeN+xxqzrLMgG5aETCBxOJSBwq63WkrrC6BdGf3YPOUH9dTnEouILLTCaEhwPkg
Us11PCyLvCtZ+yqgkcFA3+RxZMI2/ODxJTfqHBcaLIoO8E7hcWWBrhZSSkOFnBq6iQBzSO+j8iCE
x2GS+kb9cu/5KR0gW7cguEYqGhDCYudRgon12KNc4mY0k2I+3AsL88dXMgXC2aG7TlvkhWTiB0fl
Aa5TV36mG9J1dAYdYDJtEDCrbkrL+GNbwIYG1HJwSKve59xO0UFxT4ss6JlyVcQDtOXSEt+xoVCn
XZVdd2EYr17D8w53dV2ZuIGxx8EgbUQXZ6/FhmEAb7UiQRCnB+JWt2FeCo8UjqZVSpLpHhLHNsx/
NACQwoIOhKmUtv8rmq0AfLsJaHof7bQLQ5dNlrghTWELy6eP4tDuXh+VTANCWtD/BppijwSVLKYk
N/D0B19tUR0BBkuGYeJ8GrVjHT1a5L5BV5Yip1l7QmeTxXw48WfC7qrz8wEFqM/7qUQuOPOujrTk
zZ8RLjAH9BTefbViJRL03Twj3rmPYit5iLsuRkoiVaBNVkY0EL85aUTIQU4dxl2DRzV1cig6f/Wg
4Ygy+RQZ/YAb89e/8oXtppdf7ntAZuff0dSTIhtq2WrsnDx6u7NDUckt35yNver4NuV1X0JkZVWG
Mh3O0pynnRXW82M6oc7XW80znel6zvG4/AHq9mP/z/aMVj0dsv7F9RTZzle3R+yjt107GsN994uc
5bGlJ240/Jq2N+GhKy2I+yxkBmRd9RGxiG/b+KfrSGZGGC7efkDqYy6WhEqXCLvl6UgcOvkGLruD
TvO8/fbjYziSTdozcDT+JLx1bBZeed2VwdPWrORY0pI52pVZRhliDEIf8rVk3Nze+7nw3pTHRE5r
Re+2uPNOi7qVC1MVnIJixYDwk3u4RMn4MrU5w/oWxdklb4O6XjMwgJ/FJRjDpiGYbqfBbRo5016g
/t5Usu41u+ReTYhYEpRJ6RgwInXTXqNDolXZvTiyzuQBUDIHdMqHBn+A6dqkjCk496VwUArXQJXU
SdA6lkGTDOsC3bSNx6GcKHoZ7mhHXYuoU8VvwdBWUKoLy8qTm92AX2pNV0h745zQHhI+gON/l65j
lb2QHjzOO5JZR7HNkZKee7TKDQXOfSOqzi2LV/Iu3svYwf2bduIc7+QrQCOMH4qKmnNKTP0tGxPK
+IxuFiGnkSQVWj3prmATQkMn4SQ4yYAhDm76T6MEVNc+h8Ix67lz9yeHvxBtsdMhK5mtgUEkARq/
V2zPCRngJc/cjyxCzHzVaeWYcTXJJICwZyl5K3IuFxNSpEzhlYlC7y0bhEO3Pxc94fqGkgLKUeFK
MDhfeU2oFgh3UNWBX6DAkGxbkqmDShaO80JRdEsel2rYExaAQ43hqcQqSCKJne0IZj2tWm1yG+Ju
o7lMTLPjc31u+7u3uxd5pM3W6Q9lkIYmhlUFR/44lCIb1wdA7yFK1jVkdFqy3iRStmubTrkEZyUY
QDv0DGUvGj77XhSZcbLCgDxTaYns791CS8/8qa4rVQhpGWSOlqbwpz/pUPH5In9GZvsc0eN+T3Z3
OkBLcYPHLd6ZuuT2mzqbiQLIkV6DapkbQdoUliS4TIZ70v0HPqLuSujtWGNziVtVynLUgfjTy3xv
fdNSg19PjWsuLzjYipcJMQwn08q7FX3qY0y2BD3kGA0kFa6U5OcebVYKYRU/PBf+EzfW0/V8IsyU
2VZ5kRyndR9vuQWBoBNW1O7U95ryMFw0bpeJImG/0Uiy6Ic8r4CmDVd6l0veZDoFoS7MXCYmBiNu
lP/0IUhIzIr1C2hqu+xKBk4Z+dERHAPtzyyc3ig2Xbnqhr8BxvDlD84dw427Aof7IY7++FFJow5Z
qR14Mvln3zh2OpB9F5nw23coLjpuYN3Y+wmG4khwH8B6Cm65pJ5j7ezQS+zMcSIShSSeZ3HM0hkj
l/QPsm42+gJQoNeIuAK5rX3VzmZ2jlxtXM7anG8cN/kus6kyw7ih2UlbBglDSL9lai8aU0iDZeFk
OgMap9lz6lSh/Xco08XAidxa9T2KMLRpymy0qqLkpTcqcsYX0Sf3ap/KvFXaSQwhacyUk1bSZrN8
dVkpRlCmBZtgh+px2Qo3tQ/ssskVr+5oxSUpFiyeFhCqdBMduVB/XEpX3h21wRWKuBNbkUUyBOO2
qzjNkdnXoz3nz+oh58RT5D7/PHKMJrx6aiLsoJ4ktTUXI1kKOuXdX/32vU1EySJDucjXjxeHy8Gm
1EftKqUllEb0ILMETpzz8Qq8oggd579pkZaAUXwHqLFh7w6pyXMbbP78dpew/+3b5lLid0Rmln42
zahdlqYLF3zf50mv+ZKdB6g+eEQL1J83r8PJpwYorM1myxyUMgBwsuEgpX6O5SAfagr/v5OvwmZZ
7WTaLgAYZ6M9lbfLpXhnVWUkF53/49Egwk7QuwzqSpJQSgektGc58n/6QLIGBYSbPh0xa9EqvqMp
kb9C2mWUTA+PoCJPR8adKQQNWaXahdRA66swXtZURgS/26N2qpXFh5/sWo6I89AliyYydIpQnV6n
ipY3FPvkUraPgscEPCFhbPgmvIW1tNEX2bPGJiSQAYX95TCZXqOyKiHNDiW1NWz/NDd6ZthWixOn
VgPLxNyXO2XLiYT5ZlOptLpLFO4RM3XiTu9IntyMcBLcQTlzADsiZgnvEYKk4a3rrGVaIBa2U0Ct
U3zLIErduCY6b4YgH2hKh8efPmNe07ZvZkczTPir1Vw7WUrEJ4UvURRmWQ3Yjd/CTwog6CHB9hiZ
bvAUHXGyFZQLImkOPaXfJBlUv7P1+Rc7DwiHgYzZ84j3u8FFBw6xnBS/8OcTWzbH2quJPwPuUbfX
PGvsra9xYohkPjbptTCuRsE90c4Jub7gGqqcd0iwHTADipHfqgijJ4YvQ2s5Hj4Rct9+sziDs3Ve
Lwo2Wgz3Zejmye3NxZF8BypDf4doU3uHsyJ1UmpAXrTeGSoMCWyQEq25ElmABeAOTmBx/LaIYHEz
GsMc9AK0rNYqlEmiQec8XnwqCzefpS9130IyoQSY1YafeggvLb6hIMB8MB7AHLxb7/4AHBSNFi2s
+tMHlbTgyTrwpt81LMFx02MG4slhYAV1dwGjNtxMZSaakRquARCBs114TTblZyeCMPEkSEsfIS/V
FAgBfRgEjxH6Il3OUuNO8u1gsQsDognwnEZPGheumH1b/0MbeqAWbsEHmmJ75w4jFe9dN6AJLoEp
NjHepZ+KZ+Lqk5zP9FOZd3M2OmiMioVzVdsoMnzChwPdb6wDIWSog4GrsYNmbgZPhRbQxTKt1j8u
vdvAkT5907ypfG6XEdieLi79SWFQLnjJseTsXy/RYbn8zkrCndL4Tw7y77GOv2fSPS42Yy8mqyY/
c+suuwf1xaIsncqE4Y1g6m9zBje7QF0VvQF5wWMLx8Fdj74TiL+MAqxb7b71vAXuMOEe4efvmi6n
pKeSHbjyKqryaGBBkwI4uSE14oDe2+wkydpk2IK0yAWcVgviMQIFka8Je70mrKdoq9F8YbkY19an
FUCjuqg0X3oKwSPWKtGMLXtgAYIFmW1bHfeGYyYgyb4n+/g/u8Pz/z3iRsk0V8s8dR/QqWJhU7TW
e9cvNipNHRJfSne8t+nI9jGXDUAvqTiT2MtVDTsU1mLJlpSD+y4f6I3mAaSjB12z2xuT2HRg4QlV
Usprki4v9YaGScdBzir8iS1afwIKSNJMTv+RVJSh/ay+0P9iUcERaFMkF0tmwNeGku3a5BdavGH7
88Ynyg+ivc9yhV3skvsdpgplbTS031vekK7ByFXVSRlAc0lZE5qapYM0eSgwudyfQ2izvjm8NR7a
Z75pJJmcYmvJnE9jTd/mlOW7hzLPfNakpt/8BxkvnGM5O59uZmRv6Sfd1Ck5shd/9ubgR/GcMBJb
InEaq20FRDDV/49T6Mj0JvZMwh8IvaJxz8n2aQV94kpxwr6H9BVXmlDW5IFE3itJRYYzEqeN4zs3
MNDPG4ifRwtRLNUxV0kInFCit2LfBh/yOWq7a16W2nAL9nb0J6aqHL3WywKalzVa6TPta4kHM7jv
7gMExU2NsA7YChdRvWQSAWhdDNhq4gxWpISnSLheDOuuZ1M+JU1avk4sJSL9aRAC1y2nt/KBOk71
xeaxqXNR7EEp+1CTVHh3sAqGiyILo37LUx8kVv+/OWJ6KvQglumiBh1+wneRE6dDwLXxb194L1yx
dBZ49tSPf1Xbdh2M462jRo87TteJsebmlDR6YSUK94DaD+M0SqhtxY8cErMdxT3pO1AzXqELwyhO
lmVmSGwo9J9Izzpw2s68ZTKfiJ8CMFwfNqEZRjUDC5aUfK/DKqV1g/vMh2Zn1j6RWCsUW7AUQTXm
3fFvq7hCO0AdHsAJtgHBMcLCiNYBS3azp1ujbkoZLusMxepTB2UbeRY0ASYTjB+KT8c3k6hNIhik
xo+8qzD2vlbsBcDrNsDKxKihOWxC70WPtE/O4VEez26zJ1slhRJpon/mRf8lMF9HP7AAE0uT/T0x
o5dG9mFEHiISYjSq7fbukVW8FUwl5SNPQVjWiAsZBg8/ALcgpec2iP8kQg2Ri/je/LXlXvfGKG8j
8ngT5pgPxA4BpoYNuapGQl8zxm5PZNik6jRyxPxeAbr3UczZ1IscRQ0jjHJy702G20WLvTimY8vK
LSK85L5NR5wKzDKVJW29qM3kq34BurIzwNooTw4kVO21ntyx905QUDobmd0uHvNrRc+q86rMJx5c
8WmfoS/PWLkwBXILDbV/Wxs31OccrQwnjmRp1fLOAVpw0UdknN92/05SrnyYbX3Lh/FmiyCZXKub
ir5s5qFmvfdUPqRYNKMhTZhz/sZFr2JDYU9+HqFeZUAnB95tkB4ioG/mSkdQNsDyf4NllMll5Yg1
zU2hs1ZbY87Z1Ck4pQQnlTXFVFvdtytetzzU57k2ZOqpoHhqJOsV9rI/FZvr5aRWlCnuV3SSS5jj
3/zMnjbyItOoCgq138HBuLchDnc2HHNZ5LDcxqB3wkmSsihA0Je86OmyIGBzhTXjGBGEkTyeqf3a
UB/4rA4LXTMRdLTWbDOzFDnVf5AMl9AFTRN/XPllLd/KKszzQLCwyzAdXudih6p7bAHp4wcz+nIb
onwq4pzyyG8gSIrxaOzx4nMzXIZ1RKoEM/GlCX6zWWLfKEV7q6oESwMoVflHc+/ZZyVUsNZVvWya
PxKaNVwd1yk2LZIGIziQ7GZIzgQkIpcOBoTqQCc2AdnYDYNMupVuIvoqneEk5kSk5tuLZ5Zb6feq
JW9IEQ6S5Wmec4irbZ9rmImhsL3EZCymHyZk8cjJ9Eod+U/FeaGailgrYIIn8ezqyugMEXsXcEzT
/nZNoegNNL8Qjmaukt6bC1dRIe9eMghQkqigAzsawcz8rkBodWY5TU/KoXwPqWuZDP95an1ItS9B
zmEik+LGr0Y9kd1X/xUM7tPtToZksg938mAM24T7N2+CcrgkP3eT4Dh8T5i9rofi7jwozVwQ7EQ7
lUEy7Dh/T89mNjzs+pyTYPyDyX5GBE/Y66/EOpCuXIziKZ9Tq+4j3LUUU4FonTLBvdfgkOnrNhCW
MFqan+BlGv9sQBFd9yf6IA8VRRoGItsMyQdzjHvNC7zsLjVl6cF98OzJCs1a2StF2jZd+bF6orrQ
nVscehksIVY6aL/TXrHZ3g2uG8SZ5qt5ZKYAWJz1SlDJO7nAvOf5uoWmME2bxSr9rpMJPwpuw0sG
5wSt1pW0Qx7K9uuevQazRqCgqMahdRJ3Vpm2/93nYBQX/MhUmp9joEHITFU/fYg3ZmQs8GdI/uHn
8MpzZnTU5n8GZnd911l7I5s0GJQGusT7orMciBeqpX5flVhn78i79P5YW5fcIJkJp1y5niLRMumO
WoGKNdIUZ8SDjOSx50CuIX7ePf/46RI49dref9cHEtxRPOevtduUEO6zUFkr+OCV5tnSq2gb2fSq
/7FYeBGqKRW0XTgPlquQ0uWfV+LelZ5xtzbzIuCUZWSXc13NFplQwJBnpPSsIpnr+AVV400YTASc
c0wUtCV3hplK4QxbWAMJ2g+q4jqPKNwNw1XtKdtMOQKEYJj5aALUMsTN88pv1kjW+Oqf/SqLIicC
fZlC65m0foDuab66uWklQzeSjj74z8FH7Ax2ijB2wed58RiEV83Kyp2lMzjF31RcCJnev8MUBZRo
JAcRLAhUy6g8s7/PvTcixG2z+ncx5NosE1TgpJZbw4EctiWmfQV/IqSNRpa53ZPx7l5RvzxX5zbL
w/5QldbCcu53iGI4mDzQvfzYSac2+8nj0GMfZZA0v0JgJqk/usf/4sMW5K2/QMGv1ReC1WPskFV8
GTZiG1W5UjxoRuA/WqDMFGWGzBgLIARElBHhVV9INcSgifgbZYNQ6K2F3jW4GVW3jgWJQOj0nfYz
H4aE0cv6t1iIFSmEJv6Juym2KSenhJ7LrOuYOlj2TguoCeQqOJizlVchezBjsJ8Xm0rrZ19GoCTM
jBTmEiLAJQNsjR33HUPBUD7KQKYY7DOnIL6T9ymTulYGdyRqgePCZzN5Y1uUH5x9kwPvbnHGhrvH
j5WVQIcDtaUMXsmDyBDHmbRHayabgXBMP5UItOi7nGs6A0zAfAsQ52Of/hdXMtG1OWo3WTznwI5J
8zSKbZH3ZJZ/SY8K43/MgO16OUs0y2fP250k9eHmak8wxEe9EPJBEcUBytnc4p0KOzNJ2/+EVtb7
6fB4mf4UIqelhoaEa3aNpbCvd5+pYjdC2Z295OxXpAGoHhdQo0Q7NaKhYDMidCCpFSQNwkdxgG41
w/P5m+6sTE/Gca5jIDZWmRz4gJjPlseWzgDLoU56TRHhqEXSkzSEsW8Bt1ERHR+bPHURZISQ7nHq
fZRlsXW5darxZ5Xw82nKByA8PV8SR9KJWBMT/SPcrnX4nyiF7g/8ewyE+nzaM23acpbZaTTHpg61
UDodVM7WycmjX1/E6UkRVs42aqciiHbTrARKnI9zjHJqBwEJDPtaXqQIRnjuERXbDfBDBmTS6x+C
/LN64Mgbfa7w1+4sFriH3DI2ckjQ+VwsNaDpqrCdT6qeDZZxv9MAdPbtmcTTWv0yDvZiAW1RK4fY
wm5DCoWg+E6Z6SZ1rDGTPPe0M921qa/ItEvZTf1mweJ454Q+k3MAMQsfd7nuNqqwZ53mLWiDKMI/
Zy45QScBAWsmU4BqQFpq60EW8t0CBCtWoDjitt9hkfPjdwcWFIqi1AxN8nOOFiVDV19zSA/9fftC
Ivy61HFR097UpOJO067jCQhHtV2IC7EOfczcor118DpHY6RawE/vnI7jym+DO5bcG0DC1NF90RrW
NcDN7B37Kvm46d8kNu76b9bsk4Gb3xEVTPZdWHzEOqAL2abgI8KRoMT2bnrqmAnqvuotk/PYbDdm
CWOxAbeHJ3i6LNuHmYNuDNGdxLvCU1mOFMLbyS6SJGorMUEY+JiiuofFsP+hEPdJMjlBxzL7S74p
SGBY3f31C89XoJSUuZUhgB4w0/xtYgnP+LJwVgbQlXNgFkCsoUkQn7SEfELPLNkb2cBlrZvWIw5O
wKB1F3C2OES8BHLP6YnGg2en6b6acjoj21IBgP4y7aOJ1qA1d5aKIKr/h5F4b2t1sOSlz28GGg1I
bnr7UYnhboG2ulaP0/ZoreJVpJcGk0YwJ0xdQHNsMtsitjTesn3mP6X/9fsSWwHZ3ejXEe6yoNi8
bUE3sQjh1hkxByfJBdgotFIPz+06YQ/jq156/bR9JjSTctt/A70PqR5zYjYa/LC5JhxnnHqvbNhf
2klJ23pFl90RVU2ZtLMIzv3MkI4+IDFgF1Gh1D6YtCi3s6Bgy99e0oXuYuxkQgqiEf2YsTvZEcL8
bNDjvwEYO59OqlGkLsrFvYidA07XzOFcm/dgK6vaPkU8gUJ6/4zei6/W+1UZJLm3Fh/eoWg2qruM
lgG/gvAPyMJJ7u8eXMxiOpIkZn7uvl+TpVH2ctM6DXyWKUccnDInMo+3LODXck9R6puvnJ1G8g0/
zbOdRrt+m4XmYsuMFhYXYx1s0ft7o3QTbjtljWiF22WaSf2eA7GdHxuXJZgVL9aHZekvAK/nFzIQ
yxd9caGQamWFr1nIw8poAGGwEPyvuvsQ4El8p9Ne+KFZHMUtZjLQpJKFnIF2k4eFi/YaGl1n6Egm
1mtWgxEs9y7bEjDsuVDsmQ7mGi0A6AKq7VGKiaq/5ZI+sKdMkXktDJ17FZv+azHfZZLOVCxQJOFv
kOBDqG5K4Zej3pWzJX1HbezWE6dSdzNF7LgF+Oqau2zavznzVg5dWC+LH89XtWWYmSwcRqGFOJfp
gdgquCarj4gihds31xvPGqge4XSKdNMTgogF07Pe6gABkGjWeLXjY9J/OSzV1IYOjfKMaBbl49Cc
u9FFlhz0LpW8f493QNn8upvQqc8VeieeJzPq8jWOCO46SFgyKDUG3pTojbe14b7u+uQ12/BCcDqg
pR+/nVZc2diUzlqaJciZdun3tHl8aeyIHcuN/xlI618IdwtWKTy63s+/+Z92CaAFaHuqKbuHmY9/
YNI73vEP72S9T4HIvueYGANg8izWpVQ9tqcsRdPy/qltlvdrHq/ip2ktmnj/97KsLr2Ag//F/jmQ
qt5KoeyBmFmmBI0ejGuZP/+kfaOL0V0kgt5IzaU3mA4kq9rs23TKzmsrttnu6b6N+gTZuqzKSOH2
rJO+qRvIoHG+s3KSJctuTZIYCGNo13/6ElB3VL9l10ksEyLM4AiGWExMV58uGzXgfIZE+yywX2Bd
q4jy68RReAXHCNml9xmMRncnt8Dxj3+8VWfqw3tJFUJKlsiFk8PFGu7jHGWUDz+1KU5WMW3XPF09
RlTwM1fWQA5HYe4Q1e3a2FUgpWwBWFHjfCSPuy9LrIpVuJPGXdHXWohNE3F+EBhCKIecN1zKKMoa
wiFAws24Vfdg75AXFdri5jsiFBWQq1MuYGMqQIWRxD85tItzqJG7drYlGWgsBJ9E41jQTpcPGr/y
lmWl2rQDzaQ66i0H1WUmkUFyr5yvC4py0D/zylbxcrUXgex26V4CUgZy7uPri7JX5IrzhtKyzCqO
DTuGgoNX0+8IqPh7f8Uml4rwR95/lnDqPam0tgwiGeTV+PJUga79htBMGXfpJxg0t85xgYw8zkiK
h7nGMV/vWTIoY6RTW/j0uDd/xiboTKWyRIvPpG1jB6g1AJQZk278oX/nrRucWMPD2C5a9DyWlG3V
5BYYXN1YMyGF+tBjItNh8CbzBMU4Zq3g6mu1+Hr5JWtbG907S2EcSiIRX+9Tasee+vbgNr6T+uGu
qjJxX5URnrGxuDqjeV2gqu5m/Z5HwuZjSOcnZ4bbIiLKISK7Rpig+J3rzoHHK/cviqDc9irDUjGn
N3ls/A23c+pa8u7txYrCH3s9i6YkI3nTgHAdb5GvK/LjA5vLfVDpYN3ft5ReyYsX4CHSjG60JGiu
SZkfM1qqn+VvQqFXMK7zAE3zys5dnNGull3zbFJskqsMSN8g3oqPb2r1fky6P2cQQcJmEnseiCWs
nBlMj5UUxmJu79idIyzEyF4nmMbtk4fNVSgkBbRac6G6xB53K7CXvSRN9w+h17+CtuEIB95YQgC2
PRW8H+nQHqDTpPLo5yC+w3xocE/JPQb/YweYCwQ0TnQG6umojjGbh9OdIyXRZRpY6jbZW/loOfG1
MkYRa87pIue27gkUxg1/4vGPX2zT+5cfe7xW8h549zItRslUf+p4dqrvZRbt9UqJLTdEHKmP0qxP
ahqt2OYRaivS9CgNAp/mDzYOUrcJ4lawbap5Mn4nqFmGSHRJTtXJci0aVU39Oqgt4x80olVyrG3D
sDFN9xe3S6E+naoiEKTtmWfhLSXTVB3QKZ2vRpj/ny13DvpH7BtSPeqkeQZUgq9rduslUXsdH75k
UDd3lQiHtb2s3hJuC/4+EyUhAwJ7kmdmG+uJRkyrOae6ISi5VXaWzGXpXuISInGYs59a39qRUk2h
5Tt/ngM4rMVLB9RAxM0s0q9bW+9DdaA33COnT6YgBIueGTts5nTqLElK8sDocD3oUIwrhvW9SHY7
1ib8loLPQRTuChpwvXRECZI+Kt3bHD7cut5puQsJIuq7VnfI0uDOasEWlU1xZtv471zXt/3IX1YD
ykyN18kqp5e0Hih4miP16U/v3XL+egOv2PbF6V33nSz5EbVXEwoyee4leddaKw18tAlF/q0pQ0xG
6z1itPvthi6CHPn92J7EnQ4JP3b1xCJDTY9RZeAPqD+iOZkxrLVSJkYMNT+DWzyEAAiMFl1qD2tm
wEKYo4jONgLuF9Utsf4QW9Fv84ZrtkUiDDboR1EwgiwwntcmhMyue7P+Un8QW+v6JZllzJrzk+0f
aU5umi1E5Y1ol+ELlgkQSS6ORuB9AZ9sz/LSfgHtW3ZYLSp0VBneOARgtc2T9jpl65/GxXHqER4w
tcC35tpDmXTuhUUjvDCD6w7ZYZfz2LW6XRbq7xB1CAt+OYy2HywNU91AQsnvRFIY3CgcS0/zw7hD
GKFB7vNh5DbW/nz3DxIqWTV4h665jeuA8ph5SvCS6VPlOcktk0RfcHGXIS8IWzvrvXywssYFwJV4
hG1+hXlrYHlapJgoepmCWpwV5YMaxA9HBb5nMjZZy8uuK4PLn3Baclji96IOrCe2+uGQhPdNwbHO
Ig6UyZ6f1V8V/Ye66q6kxjcX5Q7nvawtSzLKc6aRgwjMM0hBJtk8sYWsgYdJnW0kjutsS5O0u/2e
/9UMXGZ4inUWamQaSa23jOBO1l3lHX0yMpvKxtO/66zn2fjrx+7WczVGIFUW4kfU0agVpHW1AFSa
Gwd0VQw7O2pgX5FK8tfefODceUyrEr165XBUqzAlbH3UG39OZnV1Y6HjGbjJgV16t1fyzS3gGy/5
7gz5yL0v1BHG7aUgdT4oOiU/ubWYS8joYLNDfAOQCQ1n7WTbiqIUSGWxlql1csA2TcltkGiNDwPp
1ely5a75FYj5VlqN12I+F88mxu4ZClqqoARGJ+6SExJFv15dPal45mYYELZTe9e2pIYc5Q19C8Zc
ULRn5G1xgddxb1TqwelMjLntD8ra3u9kEig7BOtlR+t1js+kGVXNls1AhtPlbjnRs7wdWW2f2gqM
r+g8/dgtMAZGmVHLbu7OvirMK3ulRWTCU9uIDjWul2j5OD8G+U+J9oiOn6LdTrGHCnGTxjL+wT6h
9RzDMD+3w+5JBjMydSs/PWuaLT8omLcFwGoeN/C/TaoiguadzHnS1Odywp9WHtLtyklgvpp198Ii
jtbyqx+rRKS3bTRvyThp/HEaTU+Oo5tJsxTuYbB2pQofRNaQ9fMC8r2Gz57ZeMcCop3DDr20FAvQ
/9X34Ih4cC960pfqMFG1tPLM4Atpz2YIDqQ93IDR5Pof48np4OG1my3Id4EeeXRq4uFl/gtOv/8n
9LnxuULnGmxBGGCEVy87j9UJ24cBUtam8BvKXHVBkQp/ncESZUHUrwiFxBa1UpMcj4DEoUy+AMyG
oKDUN+UIKYkzM4MjGUrPT282avkMfp8jvzJkZhAfakIzNELE0XUsrCcHaerYzZDkMzFdROZxclkx
6kwWvXxiXUBuLTxJOp/6KVAC8FVYJprJlPRFXWixdfzP6FadVVu2aTJ5BHY8blgqVrEu0/oc6PYJ
FPGxGaEO3p4QMROZFVoohMvgoQwPCgds5fzoHfbJHB6TlV4DTEasx5UR26/7VHwREKIqSnQH/sV8
yXgeOuA38nFfV41yt9Teh/THaomnrydPDIYjkP8MVZLkHVY0t4a6s4NDAJRnID2VQVRuq5jqAfIk
wgaLyIb2fcvc9oZRIrb+7ySU1LerzomG64Bb+cenI0EhLVMN5O1F7NO7IJAQme8byd3kPPCFha+S
xmDJVT2II1iBsTel+6gnkBI8JFya3IKR4dsV9Ysah2op3mlMP2YWiEGAQd8dZGKxgVlYGdzINc7X
j9QCMa8Xh7mBVCivKRKc9Vqi0wRH6VgEZklw6sDklZFNUhnHq05IIemI6ogeHCL1hY0crQKqey5F
3UNgQGmg4wvIb4tKkzbI6/PEmUkRauppILSU9Xgibv9azjfKODbRMetsXAag6Z0caqzNByKvCN97
NjfAqMB81nLOf/8UywaoQrJ6t2d0pvAuX/36tg5PsvEsdfYcbbKxYNQReYoZWadxVPTx3lKIq8d2
03NIbWiR7EnGhK2FQ72O6fB3s7YnRBUwGwdM0zHNp5wjIJY8amc04/JqMdGlt6BZUGUhK1JsUoVj
fqasAFmsrNDi+01olrk4kw21CTDNvAI8ywiff3OMBZcbZH+RpO04SWlXvC4UoIPeIh5gIofp0wA2
VOjV9EWZ7PhZ3DeCLmES9AzFHPKZ2BTXkI5s4pZbzsL+zlvM3RaCycYNEdq5aXmMuFWUwmsrF0eP
F2vyzzIr68XV2+6ijg/k2//tluJl7xTGVmmiMhyYd1Zeiwwx4IS1U/BZBKBMCctPK8PFBc1JqCCi
eiOyxmacxzUVZ+a+pZfCTlhsFmUvQouy5Xqsp3CAcLArkU7LD6P781d4/O+1/3NkvRfDbRnW9Evu
/8qFf5u7lDMhmrKyWXel2ex2QvwQgsqxrrOhRAWhMrfBH3U3O1A9xQFuSNF24L4k1ezS1JFGD+qd
Ej+TWt3KCrXrfT565XVFGZHtYsniOOH/B3A1V4Q7tztUnH2iyG9mmL/ueSSi+YUIeT0rIEIPnyyl
kLyWnz1mq5Ad+JOZY3MFY2AgdR/LzpmusrtDfU9ONAHoWrUAiCf+wOsgQE7xDKyXsrSF9jADrNnb
vYAaa1cYjYASZ68jYNlqV+0yJUpRcHEt7xPf5BbfiiuQr5O3QSv5qklF0mJYvFhKcucdsb+oFId9
9QnBz0UlxgLUSqy6BsD9ghYZ/37fHVqymMJFKq6eKRksPJ1Jy5SbgcTgCYjYSUmhU9BfsyKc493c
6IEPYtkVMpFP2Jadmm1V0KlUIar/jAXLAn0s2pH/ifP8XMiYH4NYBzc7C9cmT5ED9qoha+OQhbXs
ikp/V6hNWxaRz6puJU79q7/oYxECn3zUi4UMbkO5GQjv/R31OA2f/W4OL4tqmTRwBpO4UjX0C1T2
j+/3FEk13ZqKg46H95GK2t9qpIV/whm7fvpqZSP2/PZCsPsW/1B43+dn/UKKSuvMwudAVfGOhmlA
MZplTOPsaEHcxo6+0Ks+K1JNIYs0n6Ui4lB2jy2n17yVfiXBmV4haoAaWJBPO8sV6avARaDljpMG
aC7AzmqYUcn/sqRaql3Pz5rKuUctrTfwdevFpBBkW3n1m32C99Rr3Pb7wvJgHYe5g2vYPTz+dWHZ
+ShPGuUKyAOyh30NOIU2DwGaKDY4lSTxU4Xyc8LPOjfrqgkWfRL5y0ANvCXIevO+5YTeOlkRuK3i
4wj6JmAe/OavsC9bmKXK35+XCXFRfdk+H3fwkRaxPZuQIxy+qknopPVl0pA5TpyW6eiy/MbCj3X3
SJjzW0UpM6gkyqlw93w+SeU6dxAtRhEYiwre6EdWsG7AhiTOBTnnjN7N+UrGXW0zaIC7ouRWZKUf
BC0KHozSW7pHBKZu5KBsIYg+/AD7poK3yuW7Khj8yMsoSvY9LDwhuRmk/3iK/eY26Cjo0hiHk2lV
XpakLWwOfiC/2QZh8Ku842OwRHGCw9ZT/nWNmrIkIFY8aopNNBgWGODqilYb+4S8e0G4frQCA8SK
44Dwh1RYXEZAjlrGoQfdyDPSXsrVbvMdismjQx9G1cVuY5SFIazV82m58mzbd3sczEvVrpjVemTV
5+yizka7nCFWcewugcHoycBVz0K9TBL8FFXjPHaoRIrvhMYS1x6enWgd98Cv6KXskLAKVDvdshgb
EexYORpLPm55Gzs4Ji4FO/hM4RfDWHvidf8ndOn8Pz+QTXLRVADP4EyxyTYzTq1GkKdHjghCTkXx
Or4vMDzJRqDw2D3S8UmHJNTOnbJAA4MRMy5L+/x1vw+NpIFcOYiXOX6YFpZdBU9+lU0voz0w2e/f
pSJZjOQv1hh5xJaARgflbahdvw8nboJgqJw2Uan8dDMPXGfAbo0+XPcYd52n2c7kvG+iyf5hxZDS
9UzHCynClm6U3sEOTru/Yy/KAIja+j8PeDEvJjODw4fLqll7l50AjYC5DaDVexcxQG+zHEmCzJ3x
WiIYZbjt3ui/3Z4r/5sjdiBK/GdU1tg1eX0B9otrOtHO3paUEyDYq3L/jF47UJdr3t3ti7dBvkZH
hlSh+z6gHEV148tw9yTx+T+ZthnNtt7j/lKjt6iju0HkOpPJvb+Bfxt+4bIBtVYShg3eRqSupt3w
bHpOro3WaQx00wnwZLbbKpbt5tl0GqSGygff9IbQOUshq09Y2r7BNs6bB0ILSJ8ZMGdV8lx+kJua
72Iwv6nGo7dOoYzssldET+BlCNgfM1Px9mVQo7ZliotVLHBwbjDDYXK/5Ny323m8XJvfp6RVdWaX
It8psaoFZxSX5ExIBJgWCx9/TOPxkMR8hZHcgVChd15qyEk9DjvJXetkBJyZBJGPCr3GO+g+x525
x3rtqcTDPRJWwV2q9CByrRC2q+AecOKEpJUDPXjNYuURAITbVZE1hyqNFpN21YUF/kEiA99YndEd
lrdiL2OYC7hlcUKy1twaXLZdQpzDr2YzLC7N5eXwyQEA6BPWhcMPaiKagdLld+itnD5ugIxvpXWZ
+jwjUNk62GKphSke4F3DyDdb1vMvIRliIyeeg7xw18HXzIusSErB7tm7clohO9wXCH+T2OdRJ4OE
iNL7/VmYjAlpx3/yo2S8SzdB6vi7xLgRiLe+TtRqRKLcBogY5WYzXPfVlKj3StVQQmh619a6Yoox
SiPrNVAiC6lS/fWVXOhq8XSgvcDMqCWvC+x1trrpK1aivDMFY4plPmePRldlKZh/iWH+HUtmptwq
JRtldvHL4fqzIB0tpPqLIR/EN4kFpHjm1h0lqShD606IMPLqh7Zi2++xxXEPrqjuNN0YRwhsTGXw
oTvFEqWt69exESfLAakHYD5lCRwyXU5eN7GUPoK4c+kvTpcBsuo8VWbudpQofuty+IIBhad5Ymkf
i4YNqnWQlxc8IXlnyq08rranpKNAA2/xZQvyZ/TXBJN3FiHSt7Tt52niNJw4w+ymFnhhjl5M1Ev2
jETYCw8fnYhqtd104H3dVPxLit5nkWvwDdZe3+vCiTH2Jr2fh6g4bDX17QwEfLEr0Oq0UYNz/0yf
YWOrJB8PicxXRSWizymABAMsrfSyRT0B0Rwu5rsBXIAXPGeJasda5OpenYuWiqi53yYrz96fxjFd
Qt+6yDtoFpnB/UA7M7UbYtry1W+E6s8QXUsXZJDGuUzqqyja7+1l4Pq+Z+BhvsFQOPZMx5m4fdRC
qRzhqiigX3iNK7LChghLwTdOW1G76nJ6PxQ4LmDSVDhn84o6fAU5Ch30otxBmUi5IIhfCcklrBG1
4uwlMWW7dh1++3ru4mesoSwTfL36Qqt80d/0DStg2tqG/DLRtmKhEedBA1xkCO5rP7La4/nweh1G
PJO5rGQtC2LOVq6wyLNBEtLFfXjUSr6qgbkzLWVTmGOp/nV8JWocbOq4TJYkRtoVcyVV82vJjW1e
qJm1bbH1MfNCQxsHieKaY/CV+xFnik9cqhW3G/0CtHiSeWjswh03EyyoaY4suGpY8nIT4TL6CH+g
UcCK8sJz5W2WbEhNDd+Gdt0KBFEcmCLkSZeIZnA6j67sl35mbumNeiKyd9KYTcsqWLtGsJyjIPwH
u6akCwndT0IvaVEsuXKcqX5y3MxTe83KA2T3GzE7aKPfnJeM4Ts+u7sBCZVr9JveV939GF+2kAnL
tIjIKIBUQcV25ohKtlurTa/sn6xhqOXhPET8s5VeVHr5FC8NT47I+Dsa6hhyN8IvteOImfMqNS5p
qV/kA3I7FHBgv68+MFjJiAt/zEbVBRlGhnm3G2/xQPLfaxqq40cH8VBtj/RYZUoj+nqZ3d4t8f/j
e/bjbCLinQHl++qjU+5skqTO/Ed6BCuHqlpqAHpYno8RfHmyQvqOxS6lLPryV304SJM2JZkSj2o2
8zdcgfF/CU9YIDjP+Hc9NLzKEqzUuYD+ADlX4VgBB0r2/K/C3G7QQ3nKasj5MvED4kjR90HUnlqy
Mp+hdYActbD1txnNX38AXDgJ5YAwCqw+nJa0LvzoVudSeVjl+CZkXbhbdTkaygg/55SM4lfMWibO
d92p0aqEqkSW/sAoQjMpyzq2hKBHHg/OA/Glw5vNw3/kQT9triUnffrlBM+kGWdT/8btE/QZ4DmX
tX/o1Tj39NVSygy5X3UU+bJx6znh9QiRVeadf2beA1YuRzZnER4MtPZtJFsm1HQbhYtwWRSEdsfW
e+DWM9jmYxnWqgTCFgRndn/C6Z4UeqBgFC7MfTF1m4NOLzwRDQ+G8MKN/7b2QcB6jsZfYMN8+RdV
h7YYQn4wOxnjKZo1iIdz40aTZuTsLlBt9Fobcmj+n0boG792Uf5YtPCMFOLk6iYvT19SnusQdogf
OEcgnBTHW6uUJGOaYSYQIq0VENBkzPWAJ1h8aiFbZ5xK2oCk3q+miY0I2kGpAfXa30bAKfc3Ch6s
HYNbZBiSqYafop8E3IW9WY06iYLthVmLZIwcF/ox64MQMOuoDfuxaTykBuAelhC9Zb531b/w2Rkr
ngVuv+L+dQ+fUDdcXr5U9TMAnIrJO1v67OUVIFWY9ySNU0L7hEcEHGNIz9RoFD97ttziKcqliuVD
vQk26ELcBc5/v/17QYDzSc1uWXw0/DkD7+aHvlDMswNea38dLa1cwuGIeAavOpOkfCCoIt8enw5C
fN36qYphV3E9v+88gNhIXvgrmyFREivlDcQcFT3ibZEgndxBv+R9LGF38tedqewrHBTe0r1EhCRM
hFodt7F5U4yDOT6A59v0I27js7/aF4s2Lf0t/uIP0RojCsqY6zYjRBsYdBvb+SI57vQh3Cm+lZ19
RWcR5H/ScRdPq3wuyfmy+nHaiGiQBi4k/wKRGiFQaPZYBUeOLGE+HHzVzBh9B0IOVhR4ShO4CAaa
2ByVnL9altvjAg7typL/9i7wVhX4x+I83pm0lcCI5H414yHYVgcjrE+OHg7stdHU9ZYawgGrPCT0
ruEN3IwAdXWQuJVWoY9QxHBxOFWxHRHWUDuhz2dEUeWIXNFbYJ1E6dsu6XA0o2cCMDnSCeTXqi66
8Xz5/I7ikB55emBYrGQ8j9Y67NPhdqHUYvP6tvfvHc9wv5hVl00kfnN9FGNgjutFDNPl1HMMjk7z
supBWHp82qumZFPjgOKOOU7hFCx9mkdUKlr2/lI+XPdU7KoKUF0x1tLPiYMePVyTmtxmgOvLYyU1
vDof1Zol/QHDDikE2O8utjxTYIKc0y68pxsCBinig8QOrzMNlul+eg7N3qO2UNmNth/AKSrGevz5
Az3F6xSSQhgm7kaCwxwzvMkTpkAAAGlsYQ9sxXhIFeHQ37muBjgbx3CDlTCg4wGFt4o1lmcDCgno
7u/sZGl/Y32VSuoXvSSc+intVrwhhqs+bJY2DBSBd2M1h8BjG1uN0lNBWjI+pVHC35Eo+Du4qW0K
Y97vHUZJkmnhPHRaDWMjw0wUDLLRIyUBxgyhtVly0PN3ffyQbPhKDhD0PSZ7iCuSNSu4Wns/JRM/
3WF9ebBdfXk/rHlAa5MxbzR/3S5htJXxksF/YqC9eEcM5CoeTImCupxtswxbPTMOQLu7UDBHbH0p
Wq1SUPteYNXVSibpCtfk13NQwugqyCQiYbnTxFOeiQ1JP9C1eeAT8txSUKzu6fvajI8D+nDDAeqF
hYSUWEZJAIEyeE0ExCn6lRXP5qJ7QAHat31lg5YwfLHA6lcqW2cRciv184ZcLCI+xA3hVc6AvoLh
voqnkz3s3T5ux9Q/tdv9+dHxiw3iOeFwXjPElQGjP+CRoVpvEq1cnj0w4jq1+N6rhghJs3JAP24v
qdoKQKhnsp8O50WmQMudmJz12qVhZvINTrYMopgUXhp1EVWNQqFj8wdKmPxiA2HyuYY0BzmismBi
hsr4YVW8WsICf/Lq2gD1L3txjqrNXjYn7jVMtIsqljPWXHJwcXQbIorUw9Wz8JA+p3lgxM3FXHIS
GFlVO+AduR6VVi5nRNi4bR3fPNWgpTUvJCaYn4UEbc5BfuwDTY3mFl/xtQvMP16bam+BRyOGARYC
0Av7+mvXiBQE+8sGkuWMQ4JdmFd9sJtXUGUf4gMQwjwRfAGq/g4de41hq15gV/rJ6VcYaWs7W8qA
C3So9n1NhbGd4As18BMt566XHcVaTUSYkKdxtz6y1kJPPKgmXiaeZbJfDP+Y3NNZgqiLISxSFKA3
AKIsSGCq9k9hCNnUulLGRLH9BMhAH16PjkjPZ+SbXGFvYVva/Hkoxcznb+7gVtFeg9CuzMcJC6YS
mPPCKXjwf8fTV1jNc3YI+J/Ye95o+0GClyEwwInjzRGd6Ng0b3ieesrQSzA7zedfJDKcJB2rZjDM
CMZ8o0QI4h/j92qDH4xv8/E6VKDVmsnXnuiWv5UfPgMBVgB8JiRKJIsGOcch+oAjrUPhMG3fxzuk
F+8MZHpsdNgWniWqoPu3aR5fGSFZv0a0i/SPPSAMS3GKzXUuet5h9KNOiOVo1s5bOYeJJwCfPm3o
fe1KOv8gWbEV9zDUqo6MZKSYTShihXuo2l/NMJ7+SoU/b4BHwYuez/kMWttfuStHIIka9/NGR6Wd
E1y7KZgbUzI+GhheFtWf30Rtd4vVXUnI4dqjuPzkbIhhssgUUKJvKl+gEzbutquce7s4dY+ro1RJ
w+nYhlwoE6zqztQVzbF/sFGtL+HbkfGujHcqAHDtJzRV8WIXGTaXAYFJsHv+h0xkophxWpO5b/yd
w7X0GtcNXDxSMVAFdaiRMiRPkN0KtmKujHCcpDiFrJ58IO4ZsAotdNnFm6n9b/08GLGeR3v5K2lz
unyS6hWe8azChsXialtIlBqD2H96PbKRycrZ4vkDMzm1G3Q7wrBfCY/IGHK8msO9+eZ5qoWHYN/+
n4prAc041ekt8iBsqI6BVjGWZUNki0xl3aScajFklxhipw39k43MjKjmh4RXVpfZn4xedfsZIo/R
F8OK4Of3XymK8WLFTF3PFftIR8vFFT3YScHHJ+0T41h4VoZeLCtGeYLSQ7CviX1ViofI4VjVWRtO
JnfuyOKJDfLlsc1763yqEXK3D1dxKOwgrStJr5cylrtM0TwtyWv3MKMDEPDAdKObGVFfJkdRc3qG
wblLIZmgUY9ONJWtPJsQnPygGOLj9ek46YlEMbYKTTtc+Zb+a/u6w3uFXLhV/sfZmfxHRf5DHbNx
z6SgvqyrRfgj14NXZnNEZUamdQSUtlW4nw+/UUmpvvqp2yBM6Ygvz3btxW3hskp+SpAsmdy86tRj
h65GAyEpAKKaTRcKsn1+C4h//XBNNRoGBFyYMf6VEgpDvDM6c38Pi//yddYpnOekJQQCqbqhLhw7
LvW30ZI7vO/t1K9bPd4yZbek24AsUMVFBgj9tznvB/+06ySHqVvQ4orQeFN81OBwVLaiVzy5/acR
eky6gJ48QU5Bfjc9omM5uowimzhmpIJDo96xCUGdV+rs4ZsJQjxMfz7BojJfpVorbfuDvj1v7Hix
H5Ft47N5hNEgpBn6ijIdFcmsEHjynkQEaoQcz6lu1dEONRgVTU2F8/Ee0ROFBLjizMjpNt9XyOM1
rWuy2VomY0Y7ou7Viu+aS8DPMjsymcqwnCvnMb8FecvdqGmsqteC2ODrqL9JBaMIDguF4iCM5vSj
hkdo2+AwWSyAm6c2BO7GY5WBO9NfOaeEO2lSc8YKCJIgcpqp3HyulcWuOSUw8eIg1U6FI1L+DBgB
/P1pmbK2XZE9IhWjpcymZJ9mkfB2ViZ55dI1jVNmL4AyumbkW5ogS8Afmi+pcb8WQjd6wa8yB9B5
iUFWuNCHLTNu8lLItF1UVIMzKw6/wq6JBs/C2jvWwRQ+ITZvi1x5k3OOkk/g8cYXicwXVYIePnLl
JiGU785XldSvhrJ8Pa+2ZqcCBROCM61IabkZwRSTcdRC3Opx0UAiCh1NTEOYOXx6A2oWdYPafRjO
s5T9YNjWvAI/eg9pYYaQ1O8uooLbB5s/rXsRa7ZtPisjJ2+eE57PBAujo62ElDHBrbBkiT1Cr56q
HnpdL+nDMbNUWJXkKmIrrnnloZPyaDVLP4RuGMxEH6/xv/k2eC3WGu2Vz6OPqZ+T23ICVxXg2AY2
SUXWbDCbcqUGdbOJ1XFaGnGQWMviFvbUSph5bxCk0aTi1Y+HSajsm+pMxOIIt0PEBsEvP/Wr+qS6
Hp6TG2DSljbxEoZD3IORcK909VLDeCf4lbcFKYEABx2LB52gALcDs+UdYogvMr3OeoQI05Xwqs0A
tCSiARqIGiHbZFtgEbMVbVMiUVDD9/cFfNc1bEkDkdYtEJN3hMYEBmlxwSYfytB2mTjab+cG2MTo
EtVEwWZrK4p9K5MXnNF3DmNw0IWx5JYU1rfLhoLGPsAqJwtGLX5d4KZaV2OHRBEdDmsscbmYAZsV
u2GchrHZCppIBhsz3FrIoc42tCG9TWd4DpLFiFkx5rB0qMiAxVT7VuMaRiGFCOt71x13g+gBEKnz
Lq6z5YT+cbIb6/KaLwZGa9lII4XiLk8fJR1EAp6I6pDG/jw+RZxDIQW6GLs1gfv57xvPJ8cu8rch
A9aYgYcludmdK/C7GH4uKFuF5Fe+lfIEjDzdV9UerJ5lqquHfP6FaxZN/G75sg/twtFGovnhnrky
pOON93Np0pP/LQ3Ppv97eRUvyqNwUxupVqCO2AoDjepnbQ8r3xBEvvrfPrqCG93SZ3NR10ucUL6w
d9MziFWIscsltCjz8ikP1Mix0d8msGKec7lDNqgcu1eiWZgZELM8auPHC3/HiUzJ0IFIqp0nJyCU
urIHlAHdVfkgftdRwTHCLYk3vBUrqccro+JeRsEUiPsFF7B68QKXcvuViSCHSXfVk6iMaCbzo9GU
ouNpLeRFpykzraa+3rAkBFFkVstySME3FiZSHWqKuxAhi63b78EGdBO6GOdNoqzovSPDXKGwTpF1
evm/VIa+eZ1NnWDPeDcNPYGTzEI1aFdnlr3jV648rKjeiyx3voYVMbZfJRsHqsWwebtX19mJ/J9K
L9VGyyqqxc5lzqlndU5FVA7L1Bfus/R3xGnBT0iYLz5yBX7QNKn1sTtPbMUCHN4upi58t9O4HLpk
NEyvm6XFKb4oocPjgLBqCrAslxmTDINcUxNfwKIAxOjTpseL0GdlQPhjnW4QnUDpmeh842R2v6RY
3n+2xRNU+XIpRW83nFH794fOesl1pIg6Nz8lvvGRQBiyPsPFwkdZ9sym0lxdEif7inklH1nCL1yE
+CUQq7XjZeUTPvJGUUY51xyjXkGPpaTPMUFB2OuQ4Bh/noWK61z2G/y/Mf4Z7oO+jQGknuLk9Xhz
s9pxCuKN/mHJvYt3rMynJdZbwuVjvCwVNNRMfUG4tm6KMGb4bIPlkH8/eaDzllCEWhrr8b7oVPBL
cZg36V0pGDcEPeEOarbxlVeMia0auDsOEoWNfnyUASizN+dvG25Pfn1wh5SJEvLfKkRGDk7EFIXh
faFkgu/hODyA2vsJKVu8XJLzVQPQRp/zW4Z59msfLphMk7JpwNFXmMpq3SAaLEz740Z0pNnNij9U
WjPDQq/yw2tS6XvTtYCrbFvyktiKJtryOP9d33JKMkSnj5Ev9UxnHCJgdI09jkpD2xE8HabM3n+R
56HoCBsdVr3e8BwOYMNoao8ukoDb+R5NU+GxWI7XJZMknaip+G/Lx4WkTzA8tD8pMIQ4LiG+8OIn
KKCyP3ZcFfF8UfoMneQYVisDGrV5Z010IrBSamiGdmqgAt2CkUKKm2wGzoNP03v130s8fLIo29o7
viJ8JVvIC6wmslDuaBhJ6GU4ggcgp3p5AJCJC0wPRe/JrH7zMwSxDsNzJ2svQWbgPjTjK6Ibb/my
wbFeZVQZXZY/GOrN7vmo5Jf5GyhLcW0OxLhakfUK3HotqpbTRFvQ1RPLwHUa+XJGxdBptR+k3Gqa
r+OHvyaLsyo//BTFDI3t1TX39DcU4SjQbEvqg7uIVWRiS7eC8Xe/cqlZIZtz9R9k5ap3njUMT8lw
JLgOp6A2uORdI4+lzs/2Amn4bQH5YWQkRGej91u3JBsZxEI+b4kjTs8aGxT68sSjVHnrpAJTDDc9
8DvPnchjEz63oMHWayuu5uzYxQMZgrrgA4batZLMnK+yEI+VVkOrBD0PM4wgFy72D8f9k3VNb/0P
hOVdAllsf2CdPlcuMWVdXjzMnrwhF+x+ucSDz0hGsDr/Gpq8iSSiYhCsNRk+bVHZ03nX0V4FqmYc
gfRmVy/GjZJ2qQiuP8920Yso38cEKqJz5MrAfTjyuR0eoZR+6Oib/OcSy7T6htNINd3+mXLX8Kmu
Pp3UKzn7x3TSuZaB4YbcgWDyHjZJua+aoh1T6Pu1L0clmSrKzKrK/vG/Lc1/rdh36IeJCdroKv+k
zZtdYV+rLaaEM4LnPumXxiA2oJ8oLs9AeyppsHEaTxRhp5zl1Te2ZZ9e4skfIxL6K8zFbZfWHwpa
5ZvGgL8gLevvUBKwHp8Qir04Pj+BVxRB9YbrvEaTBnlbimwGgqOnO4T7pUBskCoiWxsjYOU1vCnb
hQd7aqpBNE7raIS3Jr2zguuVPftHsd3KwJGa1ppPdz7Raepp5RgufslHXPUQ+fZc2CyuiLUMD+P8
Z+Q5uAa2hlWB+vV2Xs0FgOdlsYTxy6nqFq+Y6yBpmsZDTsd2LTF2ga4+GIHAnSxRRPERU1ScZy3J
tuoyqdOEhwdgO+t5psgRGLYWFCDkQBTZZRkhadHd/MXJHqdLyMYfgsMD/mrbtFrDCNoU5oI0GBom
CSB00cnLURhFNuuAIWtOnQ330+EJVNggg+JS/Y5qmKIctpNolMna20u9HP8WKwTiNSTxRLtiYmdY
zG9mhPb+A5bCQoi5RHrF76LYP9fDLv9+6btdxrsZ7xjdRmGZHHS+1n5hC9oOJhbdh2IllHZszDdP
4TIr43wrKSERut33eVNilGwtGlDV9uGE6nSjHAa/6m4Dj1pQE+GXY/fCdmyLs8gDvCDw2CuXEZkq
tNKH0gvILbRNPLene2JuS9Ab7bYg/r5YIvGpzMbM986rubt474F0ZjRDBxhlIoSNQhYInD5SuTwV
jn82cgLDkJ8IxAtNaPNaJ3Ep66RUNqknfxcuVefCqcMTEXtH9yrGbatKaAfDrMuwCph6OcZG6xNt
l4ULYjhdJtFfj1Dh9k3tlpW1b5dlV1N0b/mcBx0/X8vgvXOjIyuXuMoJmDD+iUt1bT+Iv/BAzzAS
JmDLyeL4xVhfSD3D9L+AJv27DYrzDS0ifFJ2gTJ8/q28y2w9I8cND3eZ9CSnatW1Y4nPo0TTyqiz
l5n6AZJh+WYd8Fi8lcYw2MoboHtxvwbDWflzyvFeRcOEQXBi6JQNmuCgb//vRX4wpdpZvSdxkpHH
JYByhR7fw44LhJOL7q/dr6oge1NoOtHQ7wQ+DADil059KakrMI08TLlVwpmmnC79h6oQJ4hyAidy
Elu/0dMwgEUJzsV8JIsG1gSZIFUYADA+VBCx5VtcPhuuQCGOXTEGnNyPOoF4a/ZCaFSSCyf1yH52
65PKOxVmUYwiBPjl6yZDD9cTSIv98gwHg8MCdnVYRhyTp8RJVoeqNP3yK9FJ3z8q2YSs7xNLjKsd
TbA/LK4nHJfBk9dGNC9guYPxpo7tBTocjgKpRt1jIBub0V8AVrHS8TfvpIDkqZR5ENx3j0JcGAVX
VErsSSbHkswlA9Bj08GycQ2vgmqn6wwVqadgnccqiAvnradIISzQRvO7g9NxovfIihos2EQKv6Vt
aNS2ldJ77/4qe/NLDsak/otl6jyCrvCcpVXxZWLJXp06jeLaTTGpaKutjAdw8w09449AbHd29Ca2
EQUNuZoVJ6TADdFYxMtHEuafEV/qLnI2mYm1zEKyzNYn+8Z3ZMFhv4hA1IS9KXdb9Fq2osSSH0Nq
+KgQkDW3PR/h/clF//KlvwD4Be6cuqa9DPEcwXleUD9txvuO8paOEz9j/cXDPzMIqoKDAWZSTj3W
qc744PEkyqM81pOyxkur7JnrocRyirhSnzu7MQrVjXioxlWx66AE8piP81oDHilvkNSxKANwGBkJ
m9TjWrylD8eekJqiMAVeVo/OqqVc/CVrweSLHpvtAqt1iIMi1f8JauSSSV5RxV7Wymw725mbk8Ym
hIlq7gZ+aBOhsEvyhGTcbhk5ebgzLBcfGMWSKKSK4hYFm7U8mZHrQyVpctzldazC2dKYolrueIgj
Jef04dsQI38UF9tMSws3o1DZ/SF0yFxRYRZrltlFVTQl7PFvTkZJxamSLTGrToxPzkfIQaQsAo1D
Tm3fTPZlQPWCXm7C+f8bp6R1OCF+lLq+4F20Q+uzw0LNUAraqe/1OHKaK4kepGjjC5E0TalHcnwV
cXUc3/X+eBYAZUjU4MBqUk/iDUR8VA/B7xynHBRZfl4z6X3vs1uaXCD/zf84ORvXD4lF88nl9Nkv
hOio3AGxqtBga49KmLzZtq+pISS0aKQArp2egQrDxApxspvhwFLyIzJsUwm94NuDIEcw62LfQL4U
Mr2S38ET9F0vtYqGXf2XWVHw4xOWOy3+7By021bzT8rnB5KzBwrAYXhjA2WZ1HrBU+R9xK9x5nCK
Jnn2Z6YIV3yG3/xrjEKOHeBpvlIYazzBUZVtjGR0eg3dVCtLf4DVfKFH3uI9R2SJCYebrHmkcd0x
wy9wOZ0nwmQDhYaM4T2erUDPi8DsFBLsFw36JouSdBcLSLpRRHTGYr8tlEcLD0JqgqX9pb/138sy
EYsTUCSwwZXrMBYUG7tDEkhTiAh0ei0QX45jRMosbUHbuyyiP6IQtpmAahPaNeoC7Gz8wanFqGUP
sKl+UH1svtjSxCndCKG1/784e7lBVN9+H2oMqhjZR4QlfZH7vz+q1HqDqMXfBC/CPV6Cujd2WBn9
Srg8XlYo6BN2sGp7csQ8cT0aWzy/G5yFXp6nhkp+1TQDm363Fsw8L8GCvVQMHSW79X3cnCJL7nD3
WRQCY8Eg5U/yqBWw1mn9hs76HYTDPxEsK8sQbElFHnSAL2naUOfoBXFC4PtqiXRsO5qyTnl0R4oL
q/HwUevXAGlT8rpQcvBpqdaGjPcGE+PUTAYewRKI51JziYD4F6fa7ThAG+zFKdT4o3isZ7+6jAlC
iN3eoeGNiB15xwxuxpuYH634J7dpgpKAqCZoJ/Qx6rFG51KdKPVbp83IajBL6zvVgZATM3QCcpsb
1lOag500dnhJTxR6YWLUcRKrYAGtxGT9QpGttbgyThmJdCdXaOhTEyph1vSEOjrDQ+qznaRWtxXQ
wlJWYXe3h+JL4lk5LS+wA5olY9Cy3BWzTEkUswf0azw3jD3m61OlWijC6ao4ltYRndeZHqCkMzAM
/EhC+953QarI3M9NClfTLXiGT/0St/Cqv4jCb2NW3norN60jcdQ3KKQIzz52PTRAAcLupJ52Wpla
ysDzoF4AzwwZlw2U5b242FimBnOiYRHMq4sZKipoKY/r2WkekMvBqsR9D+m+zrAGNCL10t/vmLEo
najOUWF4ox3KsWnlT6lFnimKAQebcWb8tFycYo/LReo1k92PnYsuOCFqB8O0Rj407ndVk1ha+/Pq
Y4SaUr85ClNkOtspwymkAYjg0LHyT6SPFGfIZ3+kSVMFHlS0kWTqEJKCAxG15mZfeNjknSrCxcrY
GEeW9j6//WBtruRNl9abzYBrJTRB64qdVtKnii+7HKVOoPRgKLV33/r6EaKBI/8QXqMb86OUFWB1
S59FYx/Eh3K/g7S7jOZ5RKZOwIHGjVzi+qvzj7AvvVEn+S1zb851h3Nh2xlR4n8rzH7NXxIPXzOM
MZ7VhIL29CldswTjahOIKmWw4Xefp8NpbxJrRSWiAYtxzG0ilWHAQWZBSI8EeHPZhNd2RSiQ6S3/
fPNmrqjojtbwOhJza5ZTLBAJgSaXD5VAfnX1mPX919bYdjdi9IC1VPO6FzneI/DaDChYiJcwGygY
FcL0dlg5dNmuJPHRB44TIFOkTmWYUrp+l2Q6DTcppNPsO7JvQU1gXSBeFhesrSf0vT42MhBu0rhp
2oOosAhrwn3Ie7Hx2w3YMG8ovn3YSVXD/HxErxmligR9HhahooNJ+Ti9bAIOtn9SGqp0EPCKnVcd
b7uRq8iJU5Jqd/PDDt7dxnXP9xpYgQKIbz4nmX7+ww6w65E5zZto2i4xDIwAg5sRQ9ICXfJH/hmK
Wbi90tUfrB26uisptz9VnN4qJc+0RujERdNmu2t5jtvVt2sL9KktVyv+IF/Op+8999piGTgF3VH/
Q1hA4+qBWpmU1fdx2s614i6OnzHq9n+1zMw2JkkdDLiKUQrI8cYVKawVbbqJVN9LWZOHxcGy2x6u
gTJkzw8OHn9UMH0/vn1YZrluVtyry1kUR5fX67rsNONPf8saNJ/wTQAdVIOlVgczhgBpSPJjLUWj
9Z3aJEqFlVKX0zrx4Wz75uOJFOc8NM4DX9UWDxjATEIhZZe2sBYFzYiuVPOiQQv/UP0x7ZcnRXUr
tSevEB+Fu2M9qZf1f6VwRwBRMUUuWz6FioVzlRiSDHUJIb1ZMBx/Rd5izSC5KisFD3zFcLBTk+ic
iIDOVruMjwrG5+cF/mOo7Warmhqvln6KKHek35Xffol4j1Gur1AS/TtDcvpB/h33X/gDU8or8DCU
JxiybNnj3yGpNtvsa/p5+PII7v8ZTIwLyqSVD7+e+WZ9FoHHY+F2SDRAVs8uolqNkRZFB+F5Tg6X
6pVgSx+GLtktLr2tjH4F1yGfPfQs7yAxPsRRrFdDf0oUDnT63wlvaY+Tsy0vvnr1/qCDwTyePgMS
YHB8w88FDIjM33XVosot5Dg68VBOIhV2R4Y1ObMyQTtGTMQM3Kdwxko+gGAmhgmk4Y74Cma2ysyl
vJukCBkA/5p3Udfk9QLpYHcl4kM76HxmWqkAT51ppc88bkEvlEC+J3F/qOgtHyyPfMPqMl75ZI4E
5+pzz8tNNd/ZdZZPkiJqqMMPKXLPwm7cZVYUA8GkZrxr5s8QC7SMuf9GLEcuZbma7OoAv4Sx7q37
6NNChDvZN6BVh+rAui9vumRT7mv148LynmXgB1yUrp9wUKcqbZtJnuGZ9lXdR3TNxFuvXVA+8Wvp
n7opZslbEESxYdzIgX+oTHZDQ/M3J4Csc41Vnzj7OmoATodW9Tos6L7quV3VYl5w3khOTABcvJQn
B56jTThWJz9WjnvBx/ZWVxEmz1W4Z9++IFbRnRa/wFWOtT+LI4sobPOXc0bqxnkbyybwG2c6zx6m
xVKSGR/UwtLpUiIZZW1euD5YSHD1yhjYvq2jEum+GnS5qzanCFXN26zIOCE2F/sKmHQEM4JkOFha
I4TyW5vHYa17snzQD2x9kAGww8rjLG1I6e6ulaAtJl6r5HUtWzVB+OeoZoShL5tLconXrZXqksiG
RjAc7toCfnJtRqKLw+vlw5PWy54qVLdnn5gbKCYcLL/sjTW3Z7vjCaYTxcpbFMwwt16dHPKDZbnv
cZs9M/pCo+EnfA/H5KpNuxes9KHGvlKl/uqsHc0aNclBHMZCdNHxTpS1Nd88l3NRgithUjhjzJVt
1Amqg5cEfWNHteW3BfctNAG/Tltjp1gfWjK3G/CCOX8u6cl0KfHLH1vkD0df+l1gLofg1RwBbEJR
EOUMGJ/xa1wlKB7PXcljzJ+yPSfZ/UGYq6iLbvsWh8fB5EB+0z3xUadpWEJscF+deNWjBsWYSVi7
QZSTXGQI7OylbR8uN4p0BtUzwsI1oAH8t/AKttbx3k9vtsam2Y6465ZxnrKI1Oiq7vTNjvjQ8wq2
twOACUdNUTXzseT3GcN8hI3U1EDDhWvoSuBs/xMZa8507U0MkqQh8un0sEDJWxIraQtxe+wqQDYs
beFFeOaTNxgB+qxVt4bzuWJy9Fv2c/ZRKgr3yg2BZVbuFfdKtIFSGmT3FvK+kPhOmh1IadVda/5x
utwSW58jrQoO9imRJxrklX5ifnij/agVRApduF6DRHl+t25xNpnrUUZA74fM4FMl9pf9QXptHoVW
47nB4SnKPJQb7+WjElVsa555kfX+wz3xq3bcQhNY1o54cnp6RztXwEOGUw1zNlfcbHSOchIUJzLw
ZBLmYPIYxBvPZTE9wowAzB5Bqjns4CarmYefI/00DsYwDFCkrPzxHTp28scDpSZsS6hrTRdMThyV
GZlqctWL9h9iLx5wByt18pa4k1b59mr0CYzUPdznyqgaCRgcbus2G4ttGU9i3rwlv5NQVXAY5nY3
VKhOYjA2eqkRe3AjSEYEaeyMB+9b3qQo1rpR8PuKg7mK8qf4LO+EMGGrCfwZio9WgB94BVcsVI0+
2O3/uUun1NRxHK+N8cYHER6alXdt/kUKeR+rnygWz55dGgGmgBdPAoUievkXqaqRjXoEqTkiFvv6
aR9vFzovwBWWxP0oqCuS9zVEskKkNwFz+mk/Zo9vDy7xoo+QFXs5IT6/RKcerq4NxSbeGmF6ywhs
3WVDW2X9mlpS3uqDIC4PYPHp11V/Riw7pyDsS437p/UZnlqtxfi5nrFonvLUGjls9CEhnxg8uLSS
7USLjijthWRU76nkX76eZ9i9VYSGMvQfOUxexKRdrwkTLpdC9Z/cLsR0HCWHEnbesA/OhuI5n4H4
0sMjmjVUmuwpnDdw23Zw+onN//wrOHz3Qm66oxdySK/eSgYnmBAkbt+f2ESNqeNPaNZyUnid0rmV
JeiexH66Jm6/qJfZBxNOuKhcGxWGTHNorQvttirxT22Mian6y01Cp0i/Wki8DWR2gGx+qSDOPKhy
n+NL7/IfahLWazV955nbeNVIJ5tZyXrxJ2Is1AhGN3IquI8sh0LiiomZMd4/eFCpWjrC/6oVmFhl
0mfMbMBUZOaQHyzvoikdvFC1C2peTNKAd+TME3+3Ng3p02L/qYVJ5Uqcc76bpiY4WPVqtZIVeFqx
m8D6ujo/SPNl0r1AupqiTIQ/jrhUm3qHjCeCxjypfQn+TpxjI299M5K8aN0nIG9+6pzU1DByh3iW
VfjYUBmk5FXoIFlbJB0O+G3IUmOmnRqoQG97+G84dGtsgFiWcMO4hVII04T2/KJZdkJ9hfOQY5Kv
8WMp9hyw3Z5YoPwOk93kjWge2a7VIBnCLDvlMESpaq6sWf81s4ldkwNz+sEpIevwJyOiY1VKV+jP
9+OOVqsHkTRDoVcDp9b3shUoScADyPe43CecpwENAw7IDGIo9cjxYnLuC2oGT+Oiggi4AvnG+nD8
BvzAnl9k7rANyRC233y+usJYJdJ3sZ2T0Fiyl6IEYWgM818EzY0AcsKdao162DLh9OFUwIRoU8ao
uQGgKwdzC94xsjz/yD9zlIi5enpHXfhJvCYIDv68NPxSqRwubkGxhmlBFX5VNXGaWdYwD+oVygJD
6GKxb5nw36fcwUygTJotVXdxJVxdmc0oi/3Yc94edk2i0h7+l+rMs+GhNjEPc7vu12WTIYEIVThm
zCVLAwN7iECeZnHrbUhoIPMas9MuERDjFqCL9kjGytDrk6gaQzCJlEzTGWyjNmCHpvqRVK96xcQk
6UPPZynBxHpmM/1Aesy3eT2DxpACUfVfHPPhhoGGSfUtSGtPePtPAn6oJOXHJZETjc4/rfnfGOXU
MPe9HxpEYPe2OYUmkxmfvHDqb6dBgHI+LQ3LEoCxTr3a6sGh5s0rd1qAHMGSsWBV80VZDY4O/+5S
CXdnqpSDghYvemw7s9tFPcTtM+bBAEybkLCDH5zPELZgedtcYn8AEJD5ytAopnDk9R3VOOmiWYS9
UkMHjiu847vrAttRxhLkZidpeyCpqtWj55XinEYxsfQkTRJMbUec/lt8by7WvImwAGxc9RhI52zF
YSmy+dHbmDRW0RNe6t1T/c4Wa9J4ZQGxhwv3cxutS0ymGeRLxvNtQSNc9q8VnTXIuTYeQp3ZF53/
hoaeJCs051zjvrJozznLga8IU55LZWbp2o9+VneNRt3pMQX7mo2XP2x/HLsmpUh4WH36tFiHUXum
X9JIf0KtFe7RMFLiSPqu2fQ56mmlE46FzrudK74Z5MDzmz20yWnERTFfUDkXET5ZdaAWU9OTJjqP
CwTpbjFEDnr5lnU5YEO7NKFWMS8xYdSO4zs/xC0oUpr9qX7fNAnJaR5yq9c+zQZZqFWJdnm6EXny
1RynJiW+ZbX2CrLc8BqleJfgKbnlatz0xATX8F1aJYD2ewxhoy+7RB5pEv8Qttq4TbQo7SbAknk4
qmJ8xl/zbUM2a//txuEw7oVvRx4EdefODG7eu/GXXdw8/u4PzgRxARWT97wZmXMZtA31PxV89JAk
T0PavvxReOC08w8VUtHnQFMK18LJOVPxT+rt0G5cptmuYFXjKGB+adf8TuCCt/x1Ie/KB7136NJR
hJD7mUKoyCBNDR+shXfSr202yGc9h0Xoi86jLIyzDjwxLfG2jvKsB4ueoh6BRTxfRrQSLa+bkzQM
eFlYXUD0rkt6hvrCMeJtvBh1eLARZAasXZQFZMy8jzSchd6RMUax2DO/xKDlYhouKA/iHJpERZg9
trtTVUVdxgDlXP3M8xcNmXOsFGSF/Aw8HKSEenUE4LkF3qTfm5cBxlXQcLeHthHSNVjZHtxlCd0S
fV8qXO1+vUM8+SP0SIWXvZHaDQn1zwai18l5tMgK6VqfICqYiLFIFx4P4GwuxNchQXP19x6mH0so
idJ6lx+7ilvDLq7ItmCwkln6R1nDHEzCP4ouoN6kz1AOny/9+cWcBTK6MZ/a7zW/lw3JKTdmZ/fx
oNvB6HOtGGDHLPOg1p2ulqjnvcdf62+RVRzxUXZK8E0oyjeNivOS/W5GcEGuBGBD384wCZQSb9Fr
o2tE2tDD+p0pBdintKESCQ3pznWgAhXrYV41jYsdROK05NDTGKTtpjrcWw+2vN4Fu6grJ2sxrHgj
08P8MkW/JXke4dpoZTLolkMXUZyKkN0wPgliqva1Mhbv4Eb/SRpiNHYb/UFg3+O1Yj4OzXOKivVe
1QptKbOaMi6KQrNvzKCye001q23XPaOiDRe0PSs3SoVD19bfRiMcjPT8QQM3TiF517POjI2yUzP2
jFknjgKFzKpeHakHmj1YBUQDFSM4iwSALSqQu13jH+pDset19OrbJhOvngq0Hxx6mLgrPF+Dc8O0
+hBV7Ghs48/T4tgJPyte+uE6AinOSsNP6Wuqx564bkYlBsgTklGudevR/TafwUgj2aIAH49Ni8rd
hl+PTkuqQRMYAZqtMdmrL9+PnD1X5JXFdHLOxNCgtPWaxAwuFR1zjJcHUXmUcLUqkO10ZqmmYE/R
JGcrIjRC42RhpikTtSUiA2JwpmlXZvOz34gs6sP9S5GRpyttE9lnbB1Gsq0Tokl7yzqFXTYF2nQN
VpshEQnDthkTURwK4ixEJUQkpGpBKE7Bc1p96IXYW2qIOscslN+/SlpN6puBd7QyOY36D2yDqgeN
7Uu4HDKre7qBHnMk6i8p7LQmckXJ6YUr36mX+I2YDDkKqilubcQ5ft6xlrsTdiGDjEWvovzLgClt
HSvloL4YoxrNSdPeWIgN0ce3dkrvXFK3qSJgUl9Eq07MSd6gm/mi9k4PkwPODDSbCTwG8qcDgVJe
MjFkLneAWiY2HGuQTZVmnT/koj5QMBb46Z6IU0zkBtyqqE2xH0SXoMGzeqfWBXcfl7khTpf+8lbf
rbGUt+pGTF3G4qGQyGDBPY8pvHjamecHBvfr/OGBfWGJcDeWu5kh1fL7L/7pQWa9UG52ixFZXVUq
/RFu3c1pJhpIZ+6IYEzrehSQG3Vdpb7K1Q6NXdPcANBNSrV9vDX6wV6Df3R8cxAMcxmgMJZNbU4J
6E0W+5KVrjRH9zMKVwzaoDWJj8LKCijpxPguOXM7IG1Y+9keTr7CPNrYfGwmoukn1ssPFVrJAb7A
CARIqoeCQV6dpkaifyuOzoUTN92arQUTpA8v1WgT9STYOreye8OSNvZ7r8r591K5b0ggKy0P1yJh
CbloO1vU45prLM7L4CzehC0xope6uWbmtiMBzLoNtrYyt6YFl9EMhFMZj1tIOCFHEholWN1n9yv9
XGER39hVMgB7EnXjLFwVd8eMNEwvz+K3wEFh634rlDrmCJ5n6FWvhtN5U42ITJ7TdN79sbyOz0sI
EE2mLTO3BCaOmwpPzOdJ9AZbFAqUWsazoY+abF+hnfEE5fr+AMigKiIcZ2I6JAvqutI0SvvstO3T
Ah7kG8z9BH3SrQ4cxjoDRxfvs/2i276n8VdH389Dy0hjMjVQgYV992FJ1MCtcmrQg3nF2JJQZU9u
Y4a+BH6xgg6PjddTyMnkNpaqMQZF7a37z+769YuNBcBX+Nzm1UE84a3PzXJm3XhT5ACRbE+vr71o
sdsGJjDcLqEN9NeO2KMGhUYwdi0Gy/Iwi3R36A7hhuIwGhppQlU8fklOgBTZeg9Gr8ibm7BTnQ+Q
DbrcfCt4dQ0H8Z8ch5N5zoq5CNvHuW2osi2nQBdvyPJ8iyIXTHrhM0StQoCZmKE3rTIG1W4Tq0NV
f3nf3hNF2LyAQfljab94SjbKL//bqj3PQ7rhbaJCqULmyBYKstREfthfNjBgKcauCls3KghAQuwO
bnCiNUWaH3V8LRYeuoFIbRP0ikJ9xmNjfynJMdHmzt3tLxMNsOyod9DyslGwEdLxry3e2CKZbzzx
5dmW1pIsNOxfTcXD1X/v27ZbbG07ACYC+4Hv9c854pUOfBSylMqnbiID21ey96k7gtpOP+riuFLB
EzIZRcDAKCGYXGoQCyvDXq+2AFxEAmzDB7opAjguVvvQz2zfB/hqQ5GSihzJ7F+b02hwiCOZzSMB
ImxTirOSwV6EUJaTgDfmbn4EHpv78mivBW3Nm0nhPr7cabfSo9xXrANsLpGuW5dIzDDR2EWDaYNG
Th/Q6mWCXuxxNs3shjlwnfZFwk3kt8hx0aLj94G6Nb7fJzgS8yih9dt9h19QQplhVcUbE43tmf2m
yMlgrfkSkV3163I3Zuj+su8QLvtzVMOahuVNvoyvAn88lUA3tTeay6qSIpCWA41xTTs34RsVwPTh
IRqWkVbbm9z34NhwDzgXF1p1Rw2flWrT33ztW8OhXgANj5JkWtIvHE5RR7fePlZOwKGcm6jJkydJ
h65hmDDsoa5rj8MmIgRFDxllVtP39x6MPqkVRohk/A0Nn4FN4cqqa8xm29U/7mUjPsyope3sLWpU
y5xxGSMAKoIkHnqLGLp1OdI2/bbeOj50YlVXpJTk3zW5tBuVTpgK/bWrz838KTqjx+LYix0JDxy2
AZsAhEQ2nm6nqfnzObFVTXDCRNOhd/HQoxamO6QA0lytySutN/cZykoKo0Kz927kt6AnFaEsY7sa
qMaFSq223I72vX47Q0daeHbGOG3ZKq53pE/bfoGZBIe6urch+rXWY6RmJGEcbZxpnckvBpr6nkT3
oJQsEkaTRcnWKCRa4EQo/NyJTE7Qyd3m7k3Qt9iDr8YiRiqnDbIiXb2v3WfAf8CXJyw4kb9nZNh5
lg/niHYOKxGuiBhCz05djUS7D8YHz959cSEpc2tllk5B50CqesID74sZYpXBC1h9NWMtmP2v+Mg7
0sgqlnnXG0b7dAvabnp4B3Ox5c0yrtAF9FTcHOsuGQLV/brXibJda/4T8E8MjmYEagb/DadqrLyr
mZeQIVgHgKVoeeD78zfuOmfvaTFIShY335GRnl8o2ONXLm6XxRJGYpTNdE4X7RWDdz7X1kbQYwOM
0miLAxW/PYT4Ncx4OWfKOIvnzQnGH9COxrU52fCxzKISs9qSUhFO+WG1R75hxahSIR1eqKhb09DN
FRP6XlyFydHN3+alidyQOmcmGqagrUOCajTpUlzcoYvtm3/2CQ4muxIaPami5xlVo0NpnNBB1DAh
OVxVt4GPDsmXyjprE/PQtwkrrg+19OdnHrfZVFhqZLrAnpufIISgsrscvRYQ1lGw28AL3GgsJqMF
pI2TVl2NHFR7KBFdjooD+XE2yBOnjbcAJDTYIv9SaZPdrBcL4k+/19ACmziFQjKZvL2WXNk7mrvH
BXZ40uOmaK4+bkeicyUSk5/Px74SZNRwwZnLYWO7hjnnLJx/dUjs2jeTEE63Yg+z3iZhAcKHZVHC
eRs2pQB6uQ98zEsHU1f5t5XyTsWdtcWjKZRttdFB0mQ6/6DDg6KncjIrmU9zocv/KBl1Tnq75A+t
7n+KM9x69Um5KriCUNW/tQpCMfw7qoWwQg0/sxY297/9O+jnczuhi81Zy1PPR7Xs3NXnK9ORgCNz
lln0MkAG3NjelzmmCSCPwHcu2SgCAWnrModxGQkvOLgyy/Ur2v3UkUZh08u7n60lBk45dGR9hAWb
vXEGFWFI8QPcDoI2ryWuLe01JxXAGyyVZQTtB/fB7FPxL7GSw7VHFSXqfLpS5p37fTtY5aeSHqMm
ADmrzA+iVoTruoCxAJXqKCwNlHqUl2zArP3QHvrzjhAsXnqIwlw4StrZiY+VysXCjHKGJajgsUKO
d1e/wRh/cPmLFF/VBMpLPDROE53BbeOnlxEqrbUJPMprHh8peblIaIt1cMlIWfGaCkGS4vwjh+rj
OpJBkEqBA8sAw2SgSu7YkZGnZzWnGOapZow+06mOZav6xdgjARe1ptcVsg2UDUUEWXEdIRuntMBF
GkhVdPtNghDgMKg/4d0BBHlT06OfM276kcRDjDDkUBtgpiEW9mesHXF7F5yR8nIkgR0iY1xQvK5o
mo7RyAt/MM0J4VakaTZceAWN7xaqsvWZWDBYtiAGbDBRw2btDJVTBAzdEh1+xDhMrTgb45q4orIQ
yhH3lNmXxfacZafl+3JwW95NY2f5LPcRToZbTVPGu5NL61kzN9goDsZlq0vEnkBVg6IMUMpeu2Im
PvHiylJXytuG7lvJDLrkPKQrhAqCQ+kGSFqgtiFON6nqe/DeOQAFfD3aO+89SVHh8AIfH8nZQwr0
Ux6HWyt8BBxmI/QnxO1c/k7/CLC7h3vegfKyUioeUCqUETLRKqams7VXA2s/DYQ+XDJC3zeBAUEp
C21bLG9+OxauryMjOGnkqI8IJDcYc6eHL935I1i6nZhCQDjM7k3DedHTQfCcVxE/qPRhjwLxbai0
NnRpUk68v3ZCAhIaycOx43a3O9pPEfOpi87ejfBwh4YTjzw6pnqJ5DI6UYQis92Rm3y4FFEBO7L4
6f1g0MYtG7KWoG7cAeTXNGsXKuWHbuqZ8cUqezhrIDBQwFceh3pmezW0PKRvZVC3zsute7rfms73
Nfk1YhlN+4RPBMlMyCarjn8FiaqiqCE0EcbJu/cAPPGmfqStw+kULfejrKnQnAWjbULyMjpUFHDa
GiQp5NfnYk7uBb3LkjUEv/Ys9zHgh+Rj62ISOT8FnrLlP644G7r27K4PXJ4AsJ0FiTlqHZhzUHuS
6+FxFJNnmkdT+S6PRaqcE/Wz2ipANQJRkqZvBWVQqOI6fiCyn42JkmBCQY+FA5jsIZSq1eYLLwIK
dHmvmWKyXUqjPPQGHKf1nK9D29N8+Z0tiYRhuTLisWANYZPcNo1UzDEnlTKmpB3xN7fx+BnDdURw
rrAUADRuYYFqj0nGeefOry9g+WurhJCQVou9Fk7SI2KdpOmFViXo2gYoBb+aWgZhG2RsBmhMl39e
lIgkpJXSU+zF7KxHS6LXY3OTggyFagrt55BtEhyJvLxIjb66krj7Btp7bKowTB7AYzjCI4SlN7vS
SmbRifZNCcQf2xDN2IwcT5gVf2ZJPmBlgLQGqC5ARTlMpmWh2gwgLsWJP3YCa4151oCtbdP4IUeq
LpAknYo7SLkkPu9RXDtAq94L77/0qmgPlDFrz+U4lgqKdBsymu4Sejsoba7XMvOUfkJcxJhvsm2l
fGUlJX5RnmJW+RKxLkkoeNR0eW4W7Hn4XLjbhF83Z6keqEDnCH/9iNcglPNM6JiaqW0eUzhzxg1q
ssH+qYAZBJL8KBJ1TLLq4kJhY0gMjCIxRtTeuL44UM4eG6gMkraI4/nxbhOZ0N6kevhgcClCUj3f
8zWDnf/NmJ650hX392eIUZxTKbBqQcNMCSuRaI8FmGvKQCJFLpc5xO4teduTtJTg+uy3sWUWk2vQ
e44R1Emm8xj7Jn1wjfMlGfgzey6bDxkwCa8ZEb+Oap6jEvb1CP+GS0jiNS5JbJoFQpU2IMNodC0f
Zutaw6k7TfFynouhGuMb3eJ0k1VRNW3FcRgpKA2o80NlXkoSgV0nze1mOgjbFRBaCWdMhv52qYRd
TG4wsL00c4jqYkw0IrbDutbpgYwmghnbf1sy08r8tqr9c58tOmK1TnUtom6sXichs1FzeiCVUQ+T
jI7ZOiFjrf8iTgBshmrYfcDDXJHLwAvnW2ira56uEYSZ7YThikOFV5G2x1GkNk/X0lZl3RIQcM2l
g2HdcWyO7ZiIJHjZnv9pHjVobaqecr5oGcPY4DfboMkq7I7UEa9IXlJCnF4yQUz86nMG96n974b4
HgHppe0M6WlSUvL1gupmKNYStIBht8tTbOf7u1N4E+3m/DxFynqtHX8UKB5SHXadxfelWm18FBkf
1qTHy/QRapatolHUbJJsOrcCwD3jZzrbFDOOqkR9VqWz6njaN4spaVDA0OenGGGccOMSjzJJXtok
I8Di9Xqxu4V7RFvv6pzFso9W2XWsQZN2p5MCZdyR8TT5Exz6pmo6qM9BUqo2JgstLHMFpsKt49RW
rdLwprl9xBWGgYf8C77YOY4HlOYwoENj8Q4u8765g55hv5Jxz0MJatF7qiFmWxNfLnLn7bPPbmBP
DwQA7NFye7v23SBYQvTZHXqWrBJ31IoboipVwlLRFY4U6KXa49Rxlx3yfxgP0hFGlbB2mu3sGQsK
6NQJRC7E93opo5Jphjfx42kaIFW7JPSdHuA8Q5nKfEw4VQ3Mx3xK0Irk+8vO/0h2UcYLLBxNQDLm
S+uhGm1caoIgTrNG7Kz937P2OVe4jSDHGV7MSKWd6H72ayqxgN+BiqgyIJv6TRbogAfHOg12rYyB
9tMUrlg6Sujy+eO0WcbxArrJ7dpQluaQhDX7T+MZPtyK0WTD+xpV3SFNp52HF7McGlPrRU/62r0W
OZ1FoT5qbMqnxTG1VtdIpoXikK4uHXAkbWL8SE8lPrz4dwXerrfwDfn+xHI3LXleUcx+3dnH9IpZ
XDXEXVKMXsleilUXYf4jI/gzMQlFuQoJoGOJzOn9OR2rs4SFUYN+nm0scUriMjUuqiwLYiuvP2cB
VU6tvCQceQ3FEDKcvc/BZYwVE/OuujevWM8fQfBfSGUykWN5AsL7p9MKlDpS6fLvZjZGKjbb3ZvN
u195yHipa+fQQqo0teKPxSXN+75TZULVbpLCHSiVjpp2+3UC4WwR3gp845XlhtwlmXHgOAtaLaJd
ZTexZaWnOK0QWu0pOZcw4JJdlNeYg+9ih33uHbRbpl//4td9xfSFXTzSxcs+uI7yGTEEk0F4/yL/
+OBkiaGbhL+PmQkG+8rQYDpkyHJtNgtEmUL0dqUw71xlIhtYfWjN4xW36nETWoJDa6WIxWre3FRW
lY+FsIUCyFtJPpOP46E8wsXNfgF4cctWY/oLl5keKocRnzjZei86tNJ4Lx++0dalBqSM2I/tTQlP
xm1V3FCYzG+l9ypi1sfK2bj+aREW+kfIzdzsJFuic+h0pwYRVL1vijK3fyiWE+XvhhJvxvVoyLBe
ohrz78MCFlPCRdpfUUwzPV4WqDVFOk7TOwrWAv7g+fVtpF6QXC7OhhvlO9fFLHYYjG6nrMzxSxlb
Lnm08WjBsqB3rN2JcRJ/4KKeLYW40ALV6s3OTE4NxB6ArOTfYg0Hy3mpSVS4PYBEnUJfgxYGqrAw
UkXfLU2eUzFoEjqm1kQW4lubPxtng98JoYF5Lao4xO8gN3YZodiR7NzdNyBqBVP8mKQMdLtGEItX
qwL3sh+daMTPE7TLPY4Yk2KymBfsS5uzsMxxOwlybZqTKa2srEQGHY9hr+NlDEDBxZp8u/I7+W4D
VioUSoq5vSLJ/cyfae9ZPtFAz+oikXE3aeedeU7NGqy7weR4bZF0Yy4whu7IyT6BtQ72kL+O9AH8
lSt08jgRTRvIZBzlyZUHCL0Jbv/EN3l28z9Hu1+1pf9ORCET3+zL0PHE3EX+HFZuoTFnAmiIib8e
rebD8pECoO0Hpka85jfGce/+QrbdfbURvCkjHmHKf9HRp8otLL3w9eLORL3Dd8Eycx/0au16euCl
MTy//9RzWfLo+hTsGjre/sw+krXMe/vwxA5EXL+JVz+RGO5fSutglILlns/lR2ypb2yacxQR04YR
Aj7nHD2l7aBkszjRX9nz18u/lusBrCvGRFMNRXbUvuGU5dqbFyw9BRTaDBcL4Gtwv/JKbYMfRIFq
4B84bTa1bKXgxdCUgDQ5CotuexY7evndbpVXi/G4z571cT1nNj70siiFsadxSTPLLsRFShcIz16X
/3uIoqU1ROW71hutemWtsHxN1VHvPH7EMRpBFmC9ET4NQjgxdvsC+YRZMao9th3zZdOSDdTMZhN+
Mw8lvAKWFqjlZ4POnQqnKLqFQwBA+0IM61LcOT/chkwTrQwS+LK8GbWu48WjORBsvuqe2AARkc/f
xJxbS6rnXPJ4ZXAfXk9LP5h9c0OI22ZnwFAyJheKEA0MuS0Zze9859eEYIuoY2KtDOB6K5vLjGUt
2SS9h2s/6odDnT7QISDKFvn0W5Wz74sAXHLOe7Oy5E4wCH5FJZ1sxHW03VgQBSO9LQnpFy1HT9JG
3uaqoiTF1rvnDSnKdL+Alu1L4IuUij9JxHIZMyTHYI6Gf2haU6z2+xHvH0+3b6CwDT9k0S8E6Bvz
iaesigeLBYTDfADc9e0lN41QxvTmx8HA39wIi66TYkbFgOc+nh8DLG4cykNZh0XP7zg9XLsBepGb
o2fzI3qIoYWUVhap9grGfabZD4AyejQ22+svzKzWOEZPZi1rqf/pALIG+ZoTzVfGhXikPNxGqZBJ
S1uDE/o2mPAAwaBCJvEvgj8309n+/GW/5nZW7DfTmiX5rp56ZhnoShmuEtbnXsBEZQnUPr/GkYm0
0JAvoRquR9jTca2ZkdeQDWVvLvvOdSF3AG+JUlxvDXINzfgz8XqihLXtR3zvXVzTpbEdXdLWTTm1
co38f/1y8jKDt4/O1hPXVSTRb1+NuUzDGEgDIMJIjnuB3apS94RQpY6oVuGCBKfrS3vYrAcMbUhH
AT7W4l0rvXKoQ6PXzAoF5Pv3OL/sQ9FLPmfZDPASfMd9apIqPgDuY3KSaBLjzce1pprFlzmy9tnj
0p26n/hSNzTSOtsHUvJWZWU0Ly4UIr+RPl5rmiX0YjZwx11oHvNQ9NFIk6JfX7EXzp2JCMvRUTZ/
H1Rj76KvefgfDeybWiO3fTo7ztfQloZcszZeAFvoxvZ88pZff72AedQhKNCh/3rgJZGwb6Fmiyol
R2gkCTLge41Jzb79erPr3eL2vXgKhoUS8RZ8UtuPVptxkyJwmp6XQG1SBLI5MqBNd19wwmGjS4F8
XaqiDSVyFgknk8aQ8Bz4VBGTq+1X9ejdv2AeYN/MEdGOtEOEyKQN1drx86Q5jV+CdWFg4lFcjgxa
SWDEmUkK5IG7G3PbiiZDwB7T5BBVT7hRPOHKT2Q5NWgoMGoZFExhLDWHJRENt3pysfHJDABaSeBU
iNpQvPczXeT53tNX6o5P171j5OvvKVWQXHk8vrPPfiKXsfLq7HQZsHeEVxhcCWgVnRzfz3TqzZlD
pNtPlEul0pAeFE+ElQ8zMztWuNvKqfSlRBXs2/gu3Gpmb9GFYg+KD15jXfT9wx9/LzfuXlqys1pQ
HrCiJSESSmSTDXuSyD/G7Toj02B1uG6+eZmGBmHcADaaizFcDbsvnnnL26ygoUai1LBnSPSMBmAI
l5FYB+x3BCbDLIQzihC+yIKOk++tPd4q3mLgbhTTxttdDVwcSC3QjRE0Bp6CKIcCaerDV9itgkM8
cEw/Fl8wP8F9nhE3tcxa5k3ZsRcF2Qum+qbG2XoRAStCoQZvKhVaFJ/KHzn9UyGEiEQbGmKJdmHo
tM+B5i2EiYenpQQqUB3wA5wMnbmgM6bMxulkRenx2UHK8D4Tc7OlsvapWVsIgVdPKmQgxbLGJdGP
vKG/QwU47hRJBcWzpyxfk6OQmpx+XDzTwsP/L6gYj96R/c0LzlHrV9egDjR59gZmzf6pqOZBD7j0
EYzO8f16ZYVckg2Kdrr/dBqES+L5dpKrA2HyUEQzLm3Ccgn8C4vmg57CcGqw2DTPQbvS/wbmOI3t
3FyjUIOJy4WGoGNRZTZotRNg7wPjvK890Cjqu3Sebsf3yMU49yIPiprIMGESoOmJi7BciIyQAdEI
/buT+dWW8JvNvihMjz0jxNWsE5z5rzArD2ECX98PQxlRENRt3c71xNtg4VTupsOtZ/SaZln9mHx/
gsEwYQcUVABcP9gL1h3TNJZxvVOelsuhbtc3c3tdI55qR0gGlMeDEsuiqt49NghrcVmRoo6FqJhF
4NMwgsCU6VjA5Lj+6NASTSsn6f1D+INKN0UgrPNPpwSFjW9wMpp/915esuYuvgdu5V8ysz8UgvNT
/IWSI8F+uAkdt0TGykYnmVrOXBvemOMDej94PcIo3ioaAxAPhK0fVh3Q/cVjzcS/vFvmHNRcOfGy
OOziFZ+o7Cqx/YGH0JJiXYeaZRExD1Tgto0/JjtomW6wziTWtGxyTkX0LLKYRt85jvFSSLFD83vz
AiojvyeWZ5SR1owVeETHZcOydaGn4+MQvxHc27+/nRG11On9AzoXEW3n2FHEj/6HQNbHevOPPDrl
iAHMfLuMRWhVh0csyvz2NUEkHd+qGaPxrsa1l2Mt5OKDTcNQ2P3m/b88wRED9Ks6vLWN7PykRFPu
nPlXTAkOXG/F++PgeeE1IATiLITbSRKdr3XpdNmgvGb1wF3HPANNLpzHu2ksT8TZpb68RRELF6u3
y6L39vVjSHiphMOfiWhS8rqErQ7MN6MOB8VEapGggS2kKSK0m2SUn9XEfy/euwZ779BNXOpf0/Oa
frVcGPJqD00pcOJMTwu4t6v6VuajiVMfTy2vPmfaJLkZyq/qiraOlnt/jj9my0K30Vdj2Xcn2FE+
DfGZ3uE6Hw1qCSJxee+0pYofTz9uBfikQXbBzVfTldE4YFArF4mQbdu+Wc9tLbqvX/q0hCmaShjm
gdAoz3fOD8gv1m+c+z05LusPhMz4IQMDnXg0WBbfAuKODL2+6Pofh8kNtIaWlCZj3zzcmzCRv/hr
vlhmIsiiZvvjVvNXc5JMfHGIDNheHn90cUNIceM2DLro7Oa3dmL5RA3lRflqWOm4iVTQHu01WeSX
aMCFKssczcola8Uevy8G5ynwyS6+A9r/T8WGlVhswk6WGWlaFX6AMJ7344UIXn3UnuyHnJ7ZBhlO
TV0ugBZeUygITesHfkg6NaZSvtd0bcAZxidq6hREG/fnWniKk1GR5V4Jw9pZaxuelujwLxQv3uk/
rDPp9DW/TXyo9yTNUxeEUbjEiG48lEGwfhf2j4Iy8i2IOJyH1nE7DDSTg5ELx8ZcIHjaVWsw1vXq
jkeMmjUfCp9kNeEiUu4YiStwGh22krHydqyrOsGepWVOlRi4QmzOtf/MJ41qZzLdHMwvuFUvrkGu
Kt8lbbM7Y/s8rOAXvCQrM+oiu8cNY8L81K8MTIZPWf1tA5BRt0xXA5eSBa7tGCRIroV1/VkmTlmD
rLQMOfLRsI311+mdUfJP1gBqgpy5mVxejo0a13FxB8Ge7OWG/oQj+ELtvuY9Qu+elVwSoxaYCL/O
RtoJKz7odrBdk2MVi120WehaH+trqXKkR/D42Ppxz+UsOaFnXYAVwTMpb/yAvgadWLluyEAEWYtA
tK6kAu1xL8M8Fv85cn+X4i41S1XrJf4fok1krM7y8TDeLDQNytUm5OGby2s4tjdvcV7DWQxsTjJy
DUuXTeIRmWrNgEeZBEv4m7YXP+emDioguM80VS2Nr2LkjOmgxPz9e6Nfp1171xQgbtvdO0214F4u
6w6TtiuPUeJE5xbQnjvJxbz/xqpJWMVf5bQbzy9lOKOhuBugeWAvkM2skHxALccOGyGM7Th+4ZsT
brbEbeuvVpxGrukIXIqOKvirKrLfBmD7GdlLj8s1TngFaXbkXUp1DfQWOTF06zJiVuGncdjZPZBv
PWCWg4dIoExk97kklgwrreG6iTpx/ZnBjctbCTYrg//9mlQT0N8OuXVwMRoAc1hxR7hcGKPrdnGH
dHiUSNFRrTiH0FIUOKl714k7q3GZHh9g45QEY8Q4r2g4ApoJ6uW6+HVwoUzKMp+DtQIr2sRd99EL
Dmvon9eGqsuLZG2M2PEWePuMirvQy8s1vCnSzTJJhh5Mb3ccmDHuxGTd5YC9L7FtpWPMQ3hiO2mP
xhCvpXE5NTmn1IU1TmUwvx5hOo2jBM+z6RugIhDcFx0KAvZIF3UtCjIIsshLfV/yyDKgiTsRZCR0
/AcSHakyiDxCjV6Ef62Uc6lQgpYCPgn0MtaGv8bOvVLP0F7kmdcCcn79bMmDXaOpimLDUD3iW5+I
o4aIeg4kpUX45ynmYwTUWXj3y6Kfuzu9AHdb20vFdAmavW2fbmWyvKLK/FtAgzVe6YCujmH2eaUt
L0YDBP7/yCUmxFqBBucmC87NlqfVbcbLJ1QwK1n4+N9ebEU+UAB5eY5k93b3SLhl3sQf7b3bJ+c2
YzzqfY/4gfALq7Ggp/iISBpaX8DOe+LP1/N4eFznpIIUottRKUpz0QMeaM8N8yNLrvaiVoLkXBzw
VOPxRdMm243MeJ6DynKZW40jIoHP1HPGcadoxBcTQFdUyEYGz287iK87sEdijd6qJ81S5SZIgKnC
b9sHRCyrIlMg/UrZAT2TUk/enI14ppIYcuPZQQ3eRqrgK1gaaKnaa96KW/zzX1pvTC+/W58GEcnn
HPExxWHRoK6mYTZ1osto3O2ttvsc4auBYXjIgokAE97XhTk1PN6doxiJ8+0jiiTuUgC1sdM37xkD
KaTmbbwts6XTNREkD8OFDVEPlwYWAkv01Hsn6KQv1Qn84TWXRy8KPE6KbNqRqJJv0bD5Zgmglyng
fucVtMgwUjV9HoiEWd9k2HJ1Cf+tEbP6iwPVLZNO87QvGQiw2r9KrAP8X+leIqmlYK79NbJMNa/X
bhp68C/1swr8PmNLZZGiGyhHvvX56YeZ2+MrEGxBtut7fiV5bAVwd/rZPK+3GQ6fBI+Sw0STh/bj
xWcVTqZf3ExY/fFxHvQcSz5IGWJPtreCONztEqtI+vGMfwIfmdxHR6owdJcQDIkXuA6mGAmCTAEv
KdUJThbu0UWlWHkuGhkbkjHQ+Pbs9jJ+8ynXJXMnGJfmmZ414TiYbIMYc40HACIw/Spd67eNoKd1
/bli8lqL50BnBte6KnILT4gfo7dfKA7h+Ad/y4WkyaiU2bMWeMuya8M5soJHWw9MvZiwcnV1qR5L
2XnOJ3AzbcesWJ2OUwsq3r8dVVbIXTkxw54hCICm7e+sOJxg+2J0U+IY7gtsXQplXDGOUkA2gHmy
dy/vclRaL2YpmgcONE8XC7IKz/qbekXDOO0KxTKLmNIfCurUJb7JfN3MEVBaof6+zLC/RuiqdHIU
fJ1mnGDS9bq4JPQZlkylzPjoJcGLnTu13YGoiDCzoUlYgfKwU1MNAxd18I/oPfLT7RIGRpxLj5g0
nq0M+x1ckIO/W8cuC6FRTRbNog1y942KEBkhxcn0pEorRTQkiKPEN+sFWsNT3cBCCrr6KpvM7KTr
PLaJQUUlMWrlN22AIE2//qKiJWb+y2ZCx6gQt7vHKWciXIKPa4vUoMVoiCHsV7UGBCu+PRLAGDqq
Yrng/KHULePTMUrgdIii4DXT0nq6CRr+LwGYqe/JUAyAZSZNKVmX+jAodkVH76tlQ7eoFE6yUbjS
r6ohFIgiHbgfPGzbmdnhNGEupxwzqnq4M4myIpenk0Yt1bqoSMFKuaC221YM9Cg9KbFo83aI0LXn
GvIb7hsWS8MQCfkT0NjYtiYPU2YnUzkqH9CPQbvIdKr89aMMWFCstLBZeqdNf0T1GcmJJZMUw1r4
qkWG+1k7lg1tDDHqhUQjFNsnklXphizvHyDMOalsWtQkCkM1OQv58B5lEtFbu/ztoHu1htp8tt6W
+hj8vkGW5FH/BkKoKw5aZxAuA8ivTj5o1fQFNWUNMjJwzckFKLoO630YwbRsfghf8BXnqSASFobW
hqB8jldaxKyJthDTrTDbL0ORZeolSKgdmcVylVPwUXCEjhSlqGLKQdW2yEXjsXuRFQI9fX5bXrS7
Ulgn2auqNw7d6Tps98QlgRhZjLidVPCSgWAwL0C+JUM+ZqnD0iUnT/wnulF75QFPxCTt7GEXPPyO
+SmtlEB1shbVWDlzc2TYpbwHkYrcILoxIntJnq+dJrc3YOSDZvQONWxtiln78JcSrKjFwCaNDgyf
PeP9W6ZnPOruFV+20rnlC+uoHh7brPLbdksdJNKIL7PkzQwF6VP5KMuy9Zp0aHzZjjbO0BTAs6c8
lsNMgo3roPOjuYec3E8nR53y29asa6cGFAcruZ667JpvTDrm7CDLy2R6zpskxZ4OhmPjCFUpHCr2
32o4wM1mibpRh3iaBbscv0Oc5EXHApJXR1P5aOmglrK4aKsAAwSwGlMO2Lu2uiWv1Hmxr2JnxDIq
78m5UJ8SVg73yE6HTMcCznHiBKGb1KFn4cgWD8DdqS5vlOmfg7pdkhZ0l12oNpNYMX16cYdSHXLp
R+XvMkJ/49EVXepy4Nqwxff2xMm4GeB1u6TMIl4pAft3yE8vsG4eCJS2atD86JSixlz0YxBuETdX
bXV7A/M+z/+Q48ubuZJl4xIX9EWTJOfEmr2FJ1wYEpzXOu1/fOzsYmIk17BT56249spzl4TrF/h2
D9JaHxPbuLF8K7CDUO8RTzZkjRDsdj2ChPgOOnf3u1qYeHdPkhW329mVAncX5zWHPipa7Rv2BJCj
JMvUol/9DRA2QszBjB0XR9nujyhaoPjqHQYjlFmAHbycK2Qn17CpnkmSKpoYIIfiDlcX2MUCOqPW
xZ+N4jq4JNzKq5byeFm2VzePYfvMHNQvzPzmXALWNlXlgxjbthUuY+5N22PxSSV/Yq7VXjZY9Gsi
eowZb2eKesRBhaxyG/BERAmSgwIAQEty5faJf6cPOMnwU5NDapxywTayUbGx1mTpNqwsqPlKdG90
TXCC5EowtsN0t2R1aXbIsp0gAxXQ+cHPGz5iOyXQ2cDAPUuOPhYU403M4fPfvbHUCWapUqnNQWDe
1BBZPmLI4CdBtM67rKDvO8tQHwY23ggu8rHzignTS8podb921kSle1OoaaWFq3zl2HWGxKwJSUpm
scI2npmxLPRSwdOpBEby7jl855qZFZzcdqPDFaHTDRRJV+c7qo3gJmvp2C750YVLtCalFpI11TYc
sKpzSurzpxzAWOR7VRFe2O0TnnSGYJu6AW61BWWC1KLowgiG5+22tdDterQ3c35fGBisrsOG0U5d
Edqfwz60a5prt3HoCr2/8w5LpijdTMbR6geRthIWLWG1M5gqkGvwJoznaZtx2FXXpR13aCCkmJcc
dO1/XyZZzP8bUcJ0Dt2IdlJpCGh83szENDaul+ignWHAloNs2IqwQVs5+3xN3vSy3rX56ccS/jXq
Lmk3zagtVBn7ARDJLyAhr6gH9iSRQWqez67pvZSlygloPeRlHLM7ADajJgIQLn4XCOwlW3CP/bcJ
mug4iVZRdUI2Wue04mGCeZ4jrQw2VSfFKSqB1eD/vLAfTUmtcJ3OF78TZzPgg49LcuQWX5oUmGL3
iD8MFBx2SIc0MCWeS79lVPPkX52twH5JMmVGxBdVujwhaUx3OKLjbMBZxTqGAQqfyhYZbHKKGMbP
nrMjOSW6oa2WheFxgo/DItIOhihZFr8UkWL+mmlJktKyoDEOkkXI82rSY4kHdk6d9Uc2DHK7X+jE
pzU6WDPmWCgQ+BSR3Bs6ZFHUw9oEkoOhNNZx/i4dBsQEvsH0Q52eLe5wO2+gP2JLUa2LiL6h0y2s
HCc2L9in+VIJo81utFLIbeYyFIjeTpGL2UwRFT1qyCFA2q33vWIaSiWAVn3UDrjxCEgQRYIFI+7N
9mdkhtyLbdBhCtQO1OohFVm6r8wtHW4XAKK9IT6OfhFAxV/QJjwUxpNkCViDoztH5hVcUej3rGb3
Yv117eP0gNScX0292antn29uGwA65SexbB4YV+0Z+RsyOO07XFh38UvMkEvTBxM0ZVUP4u5BpndL
6gfiwBKBtN5FyLh4H2Imn4i8F399A+25Bc6HnqiSIBQMl4ZrYgvtGqFALrsOPst51R5b06LIExDR
k8DdvuyoqR/0inXWmtIwbx51Qqu2Q2kp15Ps18qLCusFuLqTsuZEdtvMT+mGvX8f4Qtfh0Dvy9kq
m5Z1bWRIyk5hBFl1vhUolBbiW8O35bw4DA3p+0X8KdHS6LIe4jcG2AbG2j8nmMq3T+NF0/6BBUlD
THGevpv5i4uCmqg1NNlBR2AmIuVs+G8DluYnuniBe2nMZ380SpUSKEWzyeIiCdUF/iVwAkVkFDjo
SidYMy56dXnMgoccBiqXWSs9SHlSBwRiO8lBQEW8VkYnx7FraffzWIFMVMjzHG6CkuVt2U2cs6oj
6xWiJ6q4y/2ayk22/6Mq6skC5c+PcyktFQuwj5oq7OAxqaJGr70+dBWutrX6HnxPfjiPR+spic3p
JoESnHPIRw+gxrnXx0wZvx3TESPScYYhC5SwlgaGWilVvjoGGkBuUPfn25u5cVITvKeHeg3idORb
NHPT/T4vNHGGdXAbsmS6t10e+PAFHW0mYdRxetC4BhvYoDA2OGW3q1hxN/Q2C4HwMhfehaQlEqp6
jK7i6p1KK9cEEvGO5bbORdPhvUByXoj9PgcXwpQYEBnvYD/8MZQNsj3Na1/cN1Sxp56AbkOCXf4g
KXbMkr65UTA6xXvve6Mi7bPve4rr21NTyAkiThWmeA44Fo5DCF1HC4Pen7qmT3MnNgRkJ79JMVwb
s5emBjS//KzW6hjnGgS5JlKJuVIcqJdQh/YcwhmcFcgDTe4VSzx+xytOtjbGjYZNwvNMPiyGU/f0
dXRALSewIinfCxseiPebJMOIT4Bu1LQEwFnhO+54rr8Kyxf4reKSqa3btC8fj6K7pYT4c5twC/mQ
iPXXJxOtFAi/JlTPuP8BIadnj5mDzWj8eDcK9k4tr1QAORYaYpWHXM48JfT5wiLJb/d8SzFnxuYM
2kHL5SlfBN4XBGrNMQ10Jt/zcoAiIgWao3IodxE9pfxn5p2TFQFWHvxHd/Nlm29grlUtJFL85LYk
qdkl3Zkow5GSeQJVIOsJvTy0IbmRwFdWXkvLk0yZIewcC/ZAp/hKX6+ocnmfbL7F3EyStu3brLc+
aOiewpwwpqQjF6hVF1pQmlfBapq48uNAX2gSLEETwU2jXgdppqxAPnnxCsKOgi+oLPJ91bXNYGKD
9zuSbZ15XO5XfNKDoL+dLU4courWL1tswnxdNxF1VvGuw4fXBL3xYF44Z4IfxTAyrLOrynygypBY
E1cNPzANe5k8bCpXJX9XOYY6ZXkVEFjaZZqmMLSZU6ondYLwGWjxZ3RM8G+6tDAoZj++lMZzYFex
ZXx68fewBV/yUoAi6MYb1Oz5CKo+kjJKXkCZ0PCERqKC4VUy2veC1PnAsQcdupIx6SFRcqbCQ2RK
jQob6tR+QBSDVXsPklGmgMbRz3z7f9tT6IBophJJPNHUuN1qBGQqQGxU1QMvhJqby/lszxo2QS4z
YYo1YGQqTMr7FuW7lyDD4T2eoXGu+h3SexSfjZJcpXrSB4i6hUXjoIiUhFDInqx8pKzfJqGle6dr
KesaqrdcR9wifbasrWGhBveaMCBwdZDzP8UhqjhjspbUpgpMdApIDwKnNbQb4TRsARoDAqV52MAo
YsDipKpWzWPEaiDO3mQpTb668l3XzU8peDSa4SFpn1cbwFXcMSJV9mgzzCYAe2BPi7gxb+cPep5E
8IEPCED5/ufQhWs9NMY8l5sqWac4Bk+XLGo6oW1OHdyax7qZjWDxD9UCqEyULFJMfaxYXwPqRtpH
9gpeS0xJohvP+OQyWTWt/wdjedMvt3eS6srz7gmdtQvTecnNl6kbydqj92jhxlxlFPkfKcziQ2/W
ziPNWXEG9oQbVDAUD78+AVyThhRCfxEuDuDVc9ZnexRMuiRwZcT8DVrMtEpMTOLAlntE7LzHa46z
w5+xPxxmlluibG0/J48qhKSoZXGRX0h86esZ1w348pvAMV0VAkJMnc/DZOXMQq1jO38LxLphmaO3
OReiBfTo2yUfVtze9g59PzWRjMTpi7fQjAQdLTSKJ3bWnXKoKHVmGrpxMKzm1tPpfhoQRc6IDyFi
0vs3dIAWz6Wv2RqAX47V1DMcnX0h3YwYdjkjCB6nifQa+AFzeeAWedQsenIS8OnXqzKxxb7VIgyN
Z2lRlBgvt/aaWSVzGiji8zvYarG2lwYBXJRC5lfteclj+lQFeF8e1cyCUdLEU8H2SXJM4dZt/uiv
lleTdYYNwgOe/uszONAvbBdA3WYHfIVzFHgmtEt05Hy97AHrJnB634ZotqdINgHoeY1KkBzRfqrt
3UxGRxL1wpf8Va6+qsPkk/Mb2qF99M/rjnjPA4PGyxCmWONDPmPemScwn+v1uV5DeZLEwUpIIL7a
cp6hrpdp7557HKBYgvoRE/6+ju2ntUXP/nG/8s2yiZcHD64gvcskbPg3d68u36vCd9AgQMFiHB/D
pZG9aIV65pjGW8Hm47hhnssG+5orEBetbRWtVclTGeoyFoX8s2BQNAdq2lfozalZ1jlRS9iNvzWX
VIRYUa/UVCpHVYceOEzuy7gjyrm8sLIxEV31O9BVQMDW9QzJNsM2RKiebYQKydTkpnGDmAb3fhO0
xLAILJyCPDht6UvQUV7TkB0hENfpPTP2MuNhFOUkZY5IYY6wi+l1r9sjxCrOQB167xmlMDjJgdka
ua645NGxP5ACyA6cTQVhg/9sVF71OxWq3ZRdGs4ptowkqflRaNbIeaDQAkj1PqRlhOoEd+/DQvVf
DVFvU+tkrUUTgpF1v6IQf2gZHXgPdDaGTGVRJL/jnXCkbJaQMs3FcQ2zKLUCprCCx1bmmmFVABD3
9x2IREX1Wl0ITFBmxTJDHBft45jkr8VPJtJXliyr17KI5VS6wymsXQu2l5rMwUG+wdAKvts5TP2H
450TYr1Hz+1KCgI7oWd4ZqKHW7Z67+Xjz2ZM7FADyv6SS9jQykvwKEmDFTwJmB7y8+5QQ9zsgZ8/
9bMMBf43q+kaYcm8icHQBaqPFmhtWrzc/Qd1ULMaT2htO+pqBTuE4nr+ZalXj/22k9GIo2eGHQC5
zfkdVZBUepxbXIGX6CyG2dEA2Yn8mA4ls9VmU2IjUVkR+JfsFcORBh0xu5mLIpC6lUk7f+Z/4MNn
MInRf5MwK0WIsl4IkPfeTuoJVh2/Pr1kYx+3foDj5P5vsGZoK+pXpdR/xg7A+shl9DYU7qvKX5WJ
ikARhRSGxF+QJZdPQzJVVrItCS7os18OA5x+VMsg4im+UwndgyqAwWjEmdhSUVMdLkwt55ZKE7Qb
dvfs/J1CdIK/6piWFYYyf68Mt6BSppWlOWvL21dIX20vC29L0aL7TzeA5CjYj07wjs+FbZA08qTP
MI44lsKp8LoicKxR4DZQGrtEls2+abJU585Afaae2x2hZueDgV3FX5zbgq0cnaf/9x0Z9sge/yiI
MUcKUAddVhmfZpvNBl7wkS9C1vf41Z0iufifkaPahRtaQyIvIsxr5mMV73V5Ojc7tuQroRtJGlU7
aiZcZsiRyqmCcedigDbowTIokHnwbv8eTh1uSOitSuDNLB7+e1FFRWXH7FjepwQx8sgC9kd1YlGm
3kQEOH2TEaVXupOsReYYs4VlBBP0sSd0ajD6w0pYnPk3w3Tmgkk4Un2QlDxaQMA8uBeFjNgAVstB
7bC9bjcD4KF8cFIkKxU6tIajsUfRsVGk5RerPiLvRjekY91Na3tlNYZtwfUrcwLsPjwgNzn55/ld
I0hCLgLnA3+yhjt/DNmsZittYwnZaIQ4YR3ZYslsxnqKXdlkv+bzyL7xjVPfuDVXBhCY0zc3Z6Ss
nkWkZK4ndLSc+8g+HiLVQtImcRNqtYH71iQwtu2eNuJ01UmGMvA1tdFVfSlAeh8Wclw/fTcWoz20
qTh9brHSNEiktopfEmBSwY4jx/fKl/3+lK3yIyg8uGnyxycR6FUR5k6hGzJ39awn1QZeTBA0/Wu5
Ofn45uzG4Ch6v4/2oBI+FqvceceaHi8nUVqDr75FnjMyM7WpzqRmstgVblunACZzfQF4p4reIBD2
X3QK52paB4VA2qsOYcUZWowgTvMB4z8EMJ8KnV7dCVBW80OD/id3nvIk4E07mod3gmiCQFzxDLAM
7PxfybEAlIx5E1LepOYt/c0S63R7nNPEv8sJFoRFAi61y0KxFgzb3yCdtx8rQWQdwTFEe1+O/O+G
qgZ9Olck8bXo2wiaglNrWq0mQ30h0ytRrPjhnwj/ODLeHb6k63ty7My8WcIIB8XGiFe5VdP9U56K
v+ID5M2M971TIIyaggBdhQQVQY8dD8+qlPDcBxL6Xzy1Jmvj3LhHSxTy4Sok+3JSYShz7sYUGLK7
kKGtN/1xZ/U4N6EebnlATxFsLXfE3V9xqMlTmW6h2dnYKFVkpb3+nHKA8xWAuNtT1uM3sF4f3FDD
R46lTskid6vdb+boaZETAGw5FPRroou1RGejBdc6aUUR2Xmnv8qZQYtq+vsabpFXbVnt6ew+swl8
sud54ahbSIu/3viswIwakGt8JU/2Z75kAGUCSCMxxYTMRUoQ7WFa5fPE0hIXJBtzJ8vzMAv98KX5
N/Rb9hg/oCkVnlXIATFINtRsZCVddxMBor/BijutAH478V1Ox6h5zw1Dkd0jhsOrYmQ5Ka3a3OPT
B16AYxyYsh1aDT3qzdsDzyDBU6cZDzWq4jFlNbO64YHExrqV2+ytEwpIdPgF8OOrXXav7kpdYRwy
JIjrQ5tBzfYlkS8TBgDmzhybXqEc0DJcC6nskocFi6/FjX9AFIJ1y2cTh2lx7wLde596pZwC99+W
rcZ7db2R295PERZ6BSr8dZevAiE8eYul+CN1l4heskffrAUy1CLURj9Dw1k4MI5952703oFrU5TV
Sfs+axLJOdEAQ8w/gyycgj6dVhiepcHYrQM0nNXF44qjaxfcEtAOzpzl+EgWYJuxnT4DLTz4EzRb
IjSgiqyZp1scTGAftO9rtx2WNjkddtRSL8Du/IMuziT38SJlxHZm8HkIiY5LGCWebrZDMHpT9AwH
x/hxBqawROvKZwdYwOiIAavYLAMJAgceGmANKTbIvePGej8RPYDtVFHsDOiPLSYrtfHRbw00V0KI
znmviufTYIN+N+2Gv/xb5k9oKAG5kuylKOiNLsF+t5+6D+JFgQp6ZlZYFpvwtqcKB9+a8UDsXQQo
SWXReYlUGvD7UXpLZSsbHFDsj2sCrvDusuRzw0xj9oauRpDVEV688t6D/J6Dhf6LxKsS3p/11qaQ
9r2w6FDYP/N/z9Q8q5mJqlm9Pt0AwVN+ABDY86pfVeST+cfJlhRAaPBeobr6GHGM1eCuPdfIy0UH
RoddKVBfaDn7BuH1FQUT3t3QG4rTZDhZxS8PODKsXY6MnkXhT1DomZY1daMZk4XgokUa7j4pt6Al
p3Jn9CyfJ9tGeHXKtLKW0ezDOcBQknYw2U8aQT905o99x1GCZTGVnK0AreEPbfnKwLQTwzczz/eY
4ydJEK//te2mtmIRzRQxN6mfqQmounDUsRFUqU/ORoNqbDHuF9ih9ygMruHgZ1BwY8bPlY5rIKcR
he3XAvvNYzYtVUlEwkXl603lL0V5Le1XUquBJVB8aQHoTl3E4gfE/xXOCdViKbI//W8dPLByERH3
B76Zlv5bOa228e7W1CmJ6NsJcNtHZrZtrjrFTFY6OOoZLV1kzYKu2geDnDF+JLTRTGHhm503/uPx
PVyCjPL5fjIdIXB0rYmeiOfM1vss5NokfYjdbzt0iDwrgUtU03UX0arXe6sza5bW7vUTM94ANnoM
kj7OxagSqnxQRGaNkGXrgNqUyIq2nnenrIHWWR2HvZKiZZ5Ja6zoGrLKTwaYaJ3trHnJcwoZYDN9
TQrgQCWaYSeQLnjMfMukmp5/sqgEesYl+PqsaOUDBQRz4YgP68lSS5NEaaQwBeSxyezTHdFLzvCA
UC0kNSFO5BfpZ2+YFkJmGcVdkwFc0LuqAv926iIZ6c9NFtoK9bNBN2b+L+uKEDL8zs6RyR05Wgqs
b8huI8GrXYZMnQG6GrGYYXhtg1vYEJNOyZHZ5YA/2xeyge/lXCAbwuFesBeIwubIkq6UTJacPmtd
Q/OlOxHwtaqXzy/0f4CO447Y3xqxP74EPBEhFFP5SKdTAeyc+itjaY7rr4LKndA4JDSSfKd/V8tV
k/lKNfsjopevSwFtGClXa/eV2ZabADC+C8q4KuVi6HZc0+yR+1jB9iNtoCrYzSIkWJW4Nj7xpm3D
kEZ7sVqiH1TD4M6DlkMMLXjtkeKAUg6EupSeLy7RtDQeWOZE9aKCYGSfysTu5Hv0cNqTHVE7eUlN
A++fbaBGuJjbRfp3OJYsXRnQehsEZsgPxRdrCHaxnldqONolVB93bRsrUx1U5hhcHn7yPGNboYSU
roe57VCUHAhhjSOhvI5KhWQK0NkvPPqlCrsPdZFP/JukGeS+55fZb7mFa0uGqU7qfEGUpJddGNDD
3tt+UKHFrcfBisyIXcpgh1CdDKsjDW4aMWp5xWj+FYfIlJvYfZ1o7a0Szt1F6lvWbp1tIfWbVwyt
WWJksnmPnk9q88cg4kTPJRlzebaGxQ9Ow7u2xjiFke5beUiVBK7AMXGUbXX/Ew3cDpBLjAD49A7c
8amHWudljqGWMeuOWJRxQeFSuge71xJqBKX4VcxJF53EesJaQpIf1U2V9ieLAdUcIdYri4s6y6Za
w+jWZwsNsOc9G1+N5IWDfpEbNRgM19fV0Y5AfZByxyf+9/aONk7uOfOWg2KO3NLeeI5FSnM93VhM
rCnUV+YQ2VVpUFfaiZHMGQoZ2cUcSpyZRrWBOmFXv7AoVQQBluDE2u6zTcBGSqSt+yZWk+COEthj
l2R8qxU4bFjuvjHISHC/0Grg1WjUaqoHXmS5+1RQfL34y4Hk++PXImsnBBCvQSAUbX6rTrVKu9Ue
R2btSFpeJ64uSI8V9V7XGP6OadhzV45AdyM2hUmEIRzPRD9mnKddhrf6y8qKyAj/pVule86ZdxZI
wIJxV/2PNMQWL0kUxbuI6n8wDvBHkhgievEdcpWPtoq6N+JXOKFRZJQ8RUCO4rFnIp040q6d5Z6s
9ZuDW/Gb87TX9b5NkshjJNwcQ2RlWk6dv9+p3xXv8kxlY9R2y4YKEdPOcYmyMnwIzLekJa7kqN8f
AzHlTlkXG9xSC8kUwHwqgAb/JM163DIvaqCFttPbysoAgBJMc0CbnePrI2eE3AjrJcyeMzbvu6Qp
ybkvJJ6ksL1SJ/vsnuVwQwx0aAlViLdcWM8VkDOhVEdGOy+ndVun2ep23QqW4IDQ3CAHxOH0PLQc
lADv9uKRSiFxjoHay/Zs/o05I/+pTF6WzFET8JwaUyzH+vzg1JISyNZV0UDrm0xF1jKU1AC83V1u
LYOAVWkywoEd33V8CYojtZzOWMjXbVTl8aJyk6M5iejpxqf3WqzJ628Ym08nP+hyAhF108BpDwNo
T4F5IWaKaFgjlpEZJ0hjXKEWRQVWiVB6xJDpCbtbMqwdy4DI8K/5nWDTrzvEylXU+JQn7W5PcCic
gN6bBQuHfXnP/i3GpOSbpLdXQSPCD3fGmfmlkJX0bjquyIifHT4p2kSD0InfWJOtlq0X31b887RJ
KDehCYlpdJH31nZgCvgijRffQDKEw/7bNRYIlLCFfgEwzIDFNYF/HPrKM1OnPJlWOhyaZJodaFsi
5qccpHBTgQsFP/k9ruRDYexNt02Q8503+Vt4E8/KUYZMHPOZY2NDQADOlxPtfn2RasvQKF4Q8XWC
J3frDF3EUfIfqjfBqsg+FeKDFcM+eoKuUzRyBPlvy+kyvSrLaQ2WrLGbe7VmOgvrdPV06XvMuLJA
+LDehN+cThUiHDIXGkBgAi1n/OXrJ5TQv1f+jbh6EC9B9HAlorlLCNh06qxV6znTrvn68MIZbu0p
3oiLWOk4Z9Z9rloyZeFIPKxueIaMvJTsUfz42/PhgEgY3gvbZk73HX3YY77ZNNtIhBA3eiPPH9Fz
Of8rMVcngvmE8AFb1w5Z7tTtFSK4HmibSAsVIy9RyQCzsdJPxi7Yii0w6E4DrZDrednc+iYDzNG+
j3dm7tU90dvxhhinKoH3utpuL/HQFyhH73/Crgs5V6SQ6uUAV0jyhPCUL+MJR+ojS0kM27a6t/u5
AZ5v7pwTflxKCwUl/2kEpAtu3wQzyB4Oa1FezTQV1NGfaxBh9QxRRdKcMalMH4rxdFhSrFGG20gT
/5lY9V70iHadH93E+EVLQ9iTioy3z7kYmVuy48IhrohVoWNYHK4EHWkYCc66h2hbh41Sp7VPs6UV
+miuu2L7JnwxO5DZ3kMeOcaEUiiQk3FXhv/sCtVVipeQESBZsZ53MJ8l8nOFJt1Ch/9Na8pXTiUd
Qu0WYjUpLE4P7402y7uVt0NkT0CLHidMgkoOgmu9jKG/V/y/mUmbCFCyLoNLMpV196BgO6HOAHeD
VHlHNA5qUm3gQQTF9Ef4IWrNTDDtBy0tmQYxEXloPRFtzakewULPZlOS0929KbJHvb5tmjL/bViN
vGvegse2gNVGVxxBoJsp9R4+LZI/Fr2nkffx54C0e3LcnAYFYTV9qhA1l5Xh2Aj765qo9jPW0cH8
W38JGHozFVnP4sMW02eN7Rli7+3UCCPHhtYmWO/BxCbKI6bPYIfZB70yup/NU0BuAL6hS967U1lU
JFLHRSc8sWB+4JSJmz9jQKh2Sdxs76jYCZrqY8J1G6uAyojdihGcps58nPhEMX7mbSpE4x7SZeaT
6Sp8Ed4zaxeTNhT2NY+yYLGl/VChzD2UsemECW9Td7WIvXm1gRi7o87xDTYr/3IXaltlXUoOABwc
fE69gOtGxalk+2WVrjjHnsfWqaxI9Sq3rd1h69ISW7Coh2hDY4mZkJTZLPLKo1R1oS4pmmxSA607
k7GG39Ok+2d6sA9fBoPIJ4kzjGsEUoEJantDoif8vdVE6Nq10JXj9nKSxWI53HTSVxvy29AsdeaX
wFKE1wu67edBRN/sq90THJYAjhdyH3t3zxlocqdg0SfXZoTcFPVedqm2llsLy3eSDoA82vfmqdI7
x+nTug6aKox9Geg3aoYr3UwSYCfNxI/04fSTBcAZLP3vHA6J2pMLcwDnUXFbZMDOuUlaNUEu205s
f3C6VRe5j98/Y6JkGs9cfesUQiKywiIGw619zcl6q91EXev4yhQP7+VhsnWgGBoeKFaw0+PVRENA
YJB3TMoxhCt9nG+Xdt7UY9TLM/UiuFgP7upYO7m+qEnyKbiTxumTQ7KbGwrC1pDtrXRfkuiC7PcC
okCG/b6oAPS+gMFE+oTM9NLtJ5v1eF96jDKSKW56StSn+7AVa4oVZ+Yx6O4aNii8DJZZRA4V+rY+
LjX8hLcTL/Dmeq5qUe/U94YnC4VdzscCBYGaoWxghO5W8xLNFhUMrX+YAxbhnDZJU6oJI/3UPXq7
pIvYQ6Mz4r2DhF86EKOWTBviGB+SpkZ2dNrMQ4Nxm+srEIp+hPtFxLK5AFJuLCSMrRGATXOdX05L
kpLScO9EAVhKK7/+9KSdKvt7F+bDfXSnYG28OieXt2TORJPgY6lZAhJ+3wfVzDYG4BbQnyaf8B4v
MjfB7fsMMV5TZBBTehgsgmYl+f5NkAQCkaeuEapKxifFshLVUTll+CCIqvMmzrD1sQ4EeJL34P1D
r7f345qplyxV9E/NIu3SwnKKQ/zakLlwPTnHLditazAT/47ZSvhreoRJhW40zVDRnooPHNQSYV1I
XUExrELtZ/EHFwFECsHpy5uIfvz3keAxSnuFjwHrowwRVKxQ6L9puSDby2NxjHHygz31II5Htzt/
nUZq0K6b1NK5niPByx1WzboQ0roMC74XEXlTB+Ol+vS1P4zFxD4eydWzHDRq/GkE8P7/Sm6otBeo
dLhGaKgl9pN9263DcOAoUtIsG/eOkdwjHK/XODcv/xh05frUPK+AMNqGo7EPTHufHUYtXRDpZJ01
nKatyBDQHZqmuF/pB5MjoKYT2z+ld41cXBDoZ/MC954nbVsCjHDUXyd04EbCZPPT99rg2TXKCkKC
w43olaISQ8T+CBVPpMHclYjAimWMoFdPvCB6MAVh7+CnX4nw+8u62NNsjLbWTezrvmZW3gfO6obO
jly1r/6XQK7V/A88gMreakjcFeC4qi5hESRe/9fEGTg7HJesEZFxfzMIk7MwpgW66gQAEGA1fRYC
BkYQITCNEK8+S4tzGHpEmWkn6ZKEHkBBPrMLxjLU/zfJglcbY7gp0EQY86dd+rUW+ST8mhHSlKWU
k+3922t741fHgQ+JC/McqUxUlor+B3KQldvsDwMoh+dGSq+P8zkVcjXuG1LHmYZzu/A7iGyFB6U7
gYsrbXG7nlWonC6bmX3vO6ZVKabBHXHI0DpxjQESisNzmNc+8Igxz7NbwfBH3hykuVDcjICjbmft
gKLu7gy87BHX6T5eTv8X+Ew3boduiWF08RtJUM804jnbPV7K0bQqh7POPlSHdMySX1q8RlzkK9Wo
w5DqHxRBFlksbWqDiby7OSaJAFQNiDaKt+hj6YrNaWwfhh9nzN5xzFzfXXRF/ashsMdLzL0VB90u
RWcKJ1gcrd0v7WVcet31hq0SM4Sdd4JANmT+5XZeRGaizShhdBUgQQjJq6bNSA8kora9kUvcVl3z
iWkM0/J4+T023fzSCd1PxcmMqnuXqFNw3HSyVT1a/W+Txy9RD1kVRsRKPEOYV8kqIqNuv+ta3Ic3
gkNGnvqICZyo2PpIKSQSVWBVx8Zm1T0E9ri7XngUbAdiAVG+VRapFB3+/UF/KKrB4QikEQNsaYXr
/lFMF4d32RSPDEkOoC3b/8C4xYZuBej+dLGDrjd4nu4K6zd6FmtmqcSvN99rTLO8z6kqj97b7w+E
onLckRhtd540yIT1GaQAQV5s5jF9nkTNFZZ+kfYuEGSVpYwdbSVIfnWnyJDC21++Px2d/itm6p6h
IpOK7GjN9+dTBILEo1SUwpUZXaOI0gm3I0KDCHH+n7cthIr1xH1d8CsIW8jtNwJiwFbO3ltjF5tB
RWPPQF2G4tDzDIM7sSFMJVozO8uM1KDIofyhveyYrwRpf6687GWNWsv0QWAKHnEVvYXok1rDKMg5
v74HVyUmAD/F/CMGnXj7TLyiVwOnyD3pYE0FkFVS3OVDBUO80l1iVQ4Hq7wIpOXhERXQZnwHL/aB
jOjqqMQqnG+4i8uyFxSSxeqConT+SV+8XFLwTda9iPdtpuZSdnpK3gnbJGsq/gqExLL20//Wely/
3awo9R7Er4sBm3bDrWk4gh9edRuhNQ9EZDy0hzX7ZWKBI7brtAEJ9VIE1/AEXbd97IUv6OAb2caz
aBeIwG7tk4831dTUpva312xpwASJU4rK6UwAEL/l10G2Z7Co/31z1joHguWZm+1MxFcp7stuO/XA
aWyAbS331ud4mT7A5DPmrtdTBtylhktwbzWBwPUPCfRwn2q00ynKuHxIQQtmqhEWDLSTx4mW+NoB
Oyf9ZpZpbIZIv1q9PxRC0Oyr+qhyflo7Q/zNdForPP1e1HGnV1TyexdEau0UehidAmdLxyqrgMCL
xTwZnJSVa4neD9ndBrl7T5gE5uEh0l4gr2Aa7QNgCFX1lYUjSsobSMWCFMNjnj19mAC30ZxjpMMJ
7A17KIP/VfEnqI+MaBBM7T82rFeocpZ73Le+A6h1eA4mP9DfWo+UF4DPjXDP+BTrUDz52ed2OHaX
gsG85/CywgVYUM+1+jOdG2MZtyjvGdUp+qN3lsV+XFgP/cZ9f3ItDv1nKgYFbpnYjPvZcvFU0Tkk
OumdUx0CQ67mip+w90qS0km4oC1iqBiwlObZqdFnS56BEBpJJO6o27SgS06m7nfbw1nRwx5/Ic79
neGotEPAMFUd0wWL9FaI8yPpNeG+arE0JHG6ag2tPXAor31aUJfsjPhZ8vel/3WyZq3+mBib4no+
83BWuDgpNkFTnOW/kVT8BlWnMlhAMRjlmGpZ+waxIYhAniwbVfyF3dSSrxEBmxVXyTZwuhhG6G+X
TJPz1V8WIseLCYt+BFlbmt/ITIs30E1+9XSiMcdC2/B67bX9oS0VDoIIos3B/wiZHK1sB4d+slOj
mqggkUE1rJXFvQzasK59aYU61WviPzxZvqeYffJWQOCgxCGztOVsdbRjz9IdqOkAC8aKfQ6sHUGe
fg0d38MjAwJFl2bFSFIEdK89A/lgh3QW0PqDRSPpgrY3Gp7SbFG/Gb2rrGkoRMaQInQidj3cG+b9
/A34O5w3dzqfY95hQEs4SWvOglmHq/MGHONa/rfLc90FtSFU6GXYMCkBr/U7MomlP3kBPPx5iNDq
kERBjbMlJVLEC9Wg165JJZdl7jAbbd0+HUKK8lqCaZOBzAgxuoVXQBwO8IL/KCk/ezGoc/kVEPN9
nKQuSSNH+WhG2FL0KSXetcs8SQPgD0vIAUlk+0T5m9Aoq6iJDZNTkT+4UPzGF+i7v1IRHbJowj4I
8h3LpEfNK1yHcaQ5DZbvPbP809HllEPoVwo4yq6a4DQumqk3qdq1Bp1awXTLzJLaQh/ZopZiPFVB
gcUTJmZoGeRdBW/qWnAyLePj6BIoSGSx+cehLM+/jtttHgNZifQRZi3qR0zZmjI2b7651O1jNSoo
pLSXSdwGoIkkeWhG4kB+9EsBEHHBRfARnNs2Ywa9uZ7sjCkNbTsXtdIHPalvtbHoKhLC00nxheVa
mAY1qlNPYORCsBYCq4dnWQbWgqjxROWovgshFLvZFcfqpO//nY7m4jzDfKxdiXgg9KNSr68YH1lK
dDesjgG9pUPTJMBeUkAyRGmaLQ6YUQ4gha/zGDovMcOPQ8oojPFBOhdnfnI1ltQmufhEOy474Ec4
5M7yOyLqCB+vthxW8J8mknAEVSfYSRlJXPfGP7Fk5eo3uHtzJI/8El2dXyEGw2LpSpvehfuMNtid
O72TUPaICTLpWwu+P4x351ZZz3W3Wze4Wapo4YAuNjJLdFd0EvESsjKcXNl5+K8Pa77jh8TTZDUT
qQVKZPuXy0mn/mo1v3bJWyMy/arc33Ozx9Jbzh7s/Ro6M7+RgqzHXgOlln4nwcAErdAV3ZHUbIy4
yBT3FDYJvq8t0zi1Jm0OAzjySxNNT+XWcfZ0anzEuzPAklp1iWiVIAUROrhcxlRngNYBGD61eS1A
47Mq+rLdSg9DfAfXOJaPGBrE64nyl5werBPRfajH4lAHGtWRptYhU5W2gLlzPgbhdNRFNNXiJPlG
un9Gq8itbFGSzYNtQaybPbyTLcKgPa2b4HqbcveA3OrHyfmWBPA3Zdt0CspUYMJXBKTRSfg6hnQm
ZRtrC4LhN5MFCVjFatz3tHJDpNspysmFQLVcmNW9dC34nrAfmVsOnLveLjlWqVx+m3ZxXCKyOiy1
o7GFTF6K4zjpVvut44pXsz4Kj8D5HgROQxKiUYE8ddBiIBHq9nAFhThiRYz3NPqYGS3rXXmoXrzA
Iqq+Ni3hh30C5Of5oPFAkEnYCjXz+11JIEXGz6zEDSgX/7ycHQSJeEFhhVpLwpwvOHRByLAkZc/i
Xx2oIz5l5iQPBMP7HOQ+DuP62y+a0xeVIWClNykvfLVIfX1yP4dIPKz5M4eDe4b2UsZ3imHqpDkb
nM7IO4K2F5OGispBuM9OErMJWgv5cez0+/2PmOY0Tib0yrKs/H306IkkOooh7fW+/hIvDSaqv2yg
0mv6EPgqy0wzra/hvUXuaOJBFHQnQuEPovK465YyovB0ZiDAv0pOJO/O73p49s94tFOAamv1SqNV
orZSMSRw0RDX44OJWe480M+Ry1U+bYVadHL9eIUugEqsOb+ZG/hAwj8ytMjQWR4p4f940XTVDM3n
+YANfkgB/Vv5g0I/xn85tO9ENukjBqIEoicnShOskYqjptOYZXZnf2RO/J/IIHaw1SxS6NVTGDCt
rdq/TBowwJCstUGBZj9IR2SWBNMLfrNnvvbN4sBftEtiHSh4gDvA/Ow9XRZhP0T56mecxPfuF9Xu
OjjVL3v7rlz354pRVMzsK7SBPHe2L23SqD+v54PXBXq/uLh0S8Fm8sbarA+B1YNNiRsHwiLv+8qq
xRlDv630sbap1Rcu37FOC9uhgFsaLMWmE9ZldeF4ZefoyLU5YoHMVA+fYgNeX2LQd5FfLH9ib76j
7r31uUI7mpT7J0jgcG5elmNefCnxkubOP6sBDeaCPHrAGSyVxM1L/YmMZ/ciOXMcAskloTMvxZO+
WR/8MhlJLHFs4E+beAgiVpVHkjywCvDPyOts7g/cF1BiZe5u7qYjAjUKtT2kwP49NiiC4F0GfLa1
xDrZKA6xQE8Zz5Wzi7tkBfbcI1FHI6QMJhNVndsgpiM6ycaFdbDAPbIZZ5/LkZ3ozNT1ej9UtHrp
kUOYTvyWKgN0fOvLwyUPbylStC2ZYIOc4Voya5G1zsdejnWVjVybXWrGv4jT4h2HzH25nxwg92GG
aSdNJi8J/sZLBJX44BHCmUtvpL3JYYLr9Cs26LbqakJU6ulPpxl+WxHSwCdJXKAwtbW+J4a5MquV
dxT13O9+PPB6H8AAhiMj3358kYfqX0c8v/kX5FqSqCxPn5XLCB0R+GpspxgUashAriKsXyLC2/F6
Jab1Ak2KFxM2d2gyQGlMAXcorjvHuR9R9T2nWP//iOlm846AmILphKV0Bv7e5zg+wyZeaTl6wQjc
CzphSdQZf/QT2I8GdKIrZIUBVBtV47U+OUbiEK/Jt3uPvq7Cg+uj+eU4aM0PNB620ZM/CjOz++uM
HxYKy6K0kU2IveZNTilqfNa74XTV5k9UzhaEN7Y9Vjq1vyooUjp8ZuEjUJ7km2r9y9O8qo89naD1
NejyygR/SVxYeJpHKLu+a0n3xCm4W2oLU4rRYABUvYC2rF33sxxyjdlw2V44ExAVRzu5r1kJ6Y5u
YSyKXYGu+qRXFCqu9XCYIiF+GnCVkG3WoGnEkT3K12tHGCCmCsvzP7orgnvMya+/c0Oy0+9MJUEQ
f13eSnj1OFSAy/en+UP+0FJMLDmXVESaK0//ZKkqJv7/lksgq/TT7j+v1DVhPhri0UKUS9igI/JC
vIe3mziRYaDKs++FAYm4kucrsfn19+6w99g1dCLSgC7kE1gXv1vbyPqPhlxZZudxt+noA3RaD2lu
CKUaq4j7xSSn9tfEIB7lBPeSOJmHvXm+HuIK9PmDNrpAj4WIueCSgjJb9bSjqa/Ts7UzMZ5RuzIZ
d2aOmYh24DiC1I9lgjdxkx96wzfj/spHn7q4kEPeXPGDkmgHgJdRkApfLizqy9LLFwolAj2ltp7y
K6r3FOfHCftqgmZdlh4savAT47kSUv41WPsM6mtBaUGbpPx2gbUlmwMVXczzLnPsmOobfYHJZPb7
PNdn0gUz1v87mmt/f07+muOT7eoy8Zyw78ivIhUbwWzAuvYjBBFyec8cnlwVd0J505Zpup0323o5
jBSJe5W7eF2W9hPFEYD5A6qfSkjicgB2xuRTSkPH2JRMLRwN3II7K6o9kU+95BdL5+W61Vs/qog4
9eSCDVbiQoKO8+Aeo3XnabASIByvUMD5PUcyzx1rFeFV7aHRaCiHZuZhlQLzrRKg82+ZHOJO1M79
QCLYjpjvgGcY4n8594pd+ZQW3mZVptrGFxu1j5csKifVLqtbNdVbrRIp3hiL55sqYoe276hdcCGv
BInw7Nf3eIWMwIJ+M8USekhztOdEtSbAk0HWz+NnGHNCNjsgO+1hwfLehWyec6oko8M2MCfZbMey
JZHOFoRR/+EUO68EZ03OTiOprMd0hQrs4o/rbSFOhuTP50V7a0rlRtEOqad4/HHDM8w/4/E0BzEq
xnRNcJgsIU+8yU+D9FQ//oGTKQ5hj0I3Bogbio/Wb0rIe6B+eqFx3HAEXlOeLEQft5lGd/J4Tk4h
jg6pKmTN8PlcdvJ6LbsXy6Quc1F7oXT+oq8odzNY1sh2XR3dV1JGgzyIZQlxcDWFHuFsP/N5sDTz
CTqjnsmUZkR+pWqWR6IsyY6jfduTD+qeB0Q6wMTAidGYSfPMvYqSSvtqgrWWiHcSg/J2D1rIrwYE
LWkTdbFaVX32b/Q3PSDiev/TFE4x3yQSkSnX9sFKNKG5VX5jiMNdIT0bII9ogsXl4wtoFLv6mMnv
Ldt0BA7LHBIiSNO6Vu5/8TMV2TYbezwfG/RhvoEJwVYH+23ZesoGR+buj4i3Tw5jH76pGxtS58Tv
yDX93zDgh0LXZyvLsgEW/26WdczZxn4A2oHp0movwe3rbPIDrZtxW/3PqzxY8jHqPu+44JGX/nT6
JLR43m+dTlUIH6jkkMmLDPwhZzPAoeAazBMu7c+ZLSLviDUfYltu0eHepBcyt9MQ/7u+YM2isRSx
36mTEqjePPLnzkvMOn2VGBRYCCU7/eL8LADqelm0LgcfS9lvyNtojPm2QVnjO3u/4Y6b7PZ2ENaW
RqPRfimq6PIaqGjJm+9nVVvrSNZZZfNZQijDLmkVUqRqdcFzHSQAZgrvXvuAMaDwnLSznB4/JQw1
DsxRLbTzs2JoRhNIp5+sntJhtXcpphdFBpWODi3ozFgU0h49eAL9ck6y1/TNEpXZNnbEKy7A7DAN
45bla0uLEgm6CmOgfpF8sDiELA9AowS0RoocMBgzrDA0Dut6W/ZA6hukSF6hUb5K/QDg3CtIHaXJ
49RSqXsNuPNDPK7DxfFv2eg4diHBgPW5ELKcmv0bCPP+KHSHyPiBjkRXznvDrn8enYPZvHokYvQT
QvcsjxJuIrNpn7e/hLNpYk7eJVJPI06Zv7ookTg+Qdy53iPE4IwwASCcytk7fiM+DcuRJUuvToEJ
14Wr62m0UqIcIvDARTfGoExyjK31PVDIT0m4TvxBrPn0LMxwbkQFte31Hz4fNinVAWDYTEQBlgrg
AKG2CNYRUB1WP3myq6HcJaIglVB9x4VHyJeCUNdCJSOgupyfT09F1jtBtYr+qgqk/iUNpRgTzvje
JNbEJNgukubFLu99a99sqsqgkV8xZ7SIJc2QaLtsE6MPIIE2cWal0b7IF9UnMCR5TLmW3N0KDsQp
NTlvgbG1ekXdDTE11tYxU0MSpWkEalnLwubH5jC7mzzfKuWrt8FeKDHFRtbUEqbCvqI4Yhue0WoL
kzT7LwWJnd5PyO3xm9OVJ2wwtLFkLKpIlhnwbdCM8IUZjJgePHFtaXj0VULeSGUd2Fh/5GuWkYVc
is7aGdJMuHCwe2iFanUqa6anbW8yZG+pYnxZkkXYy8Zn0nFPlUNviHAN/bCcgB8trrSXBRuAD2zd
BTidZs83as8SuqVdJ2mQEbEN7fTy8ukcijnSXLeSBwBEF/mSkp+MH85oiuW6HYuDInM+ghG2Cg+T
U52QZBZJSXxiAAhc0SDk/5TOmzcJRrN8PNrE7nUEPVMzsWrZjTwa6kKBV3o5mIyYN8bBr5RGg+Mx
36q4tbQu3/Pjh7RnRJm3gItxyGQY8U8ro6MkDyrvVBhdI+G/Xwr8R/zYO3+QJ3V3RlD7lQ2l6fIN
uWddSZcPFuhbk8VqDKCTS0YRGGRASUEdIedz/tR1m3+tVzJNZziSE8UAdo1NSbSh4n2xCGWohJqI
5oGdRQvA78jwWfIxNwmrLTcwX/PXyuvEJ6IF0y4VLgjSLiwBnQHN7+91AxqhD9oYhddJfTJYeNVs
WUY6VSL4wJXVK2i7DUm7OyIYLdt8iC+o+sOu9Oe83od/tBSEk0iBtRiSWp6lHxAuzDf61udMrXvz
2F5cEPwziRHCEJb3Fa6T2hUzoA21gKdrlBDZKGGHuKALZqYKeMT/i9ODhz4YAFIe19NYHLIshU5t
cCTCK8pgmaWuPIwGmMOT1c7FvoclIY70ey0t5tAGQ8Rnuv6cSUplQROWcykL8CQ1tZs/Ln8GQDKI
5D/Z5w6TRMWnynZnHBd6SWcNDu9OIn/rl8SK0RoqZsiIHO2Ya3LyXgKE4pHZXkaGsGkkAMbi2EbM
6QKDOtetH0q3WNiSMBNmd3fh5b2WLO4gteIG4B0THu8quvdWci4eCpDQsaSo67gJw0QrhblphyhJ
HlCRjTZqoQtExRzi8HpL4/VEQz2nMcYSWdQq/m3VHuxs1dKbEvJ+cUNBBqquR9HBWNrc4/YUI8ei
QRV1vBuEKkvUT0CesB0iRJeDUjFOGsqh/SWn6lei4WYt9vxXj8jEm1jyhHNim4AsGbCU2LFEbCuu
9iUgKKFsNYtNfDa+in3uVCMkPRqYm2Md6jFCHysgKLv9c4nXEGV0euzOktLrSMGkb44CSucIbNpt
YLGOq70336tpECBd8sv/WNJ7RXrTQ77zsOkHXgvrjkSyjy1ONSy/2ZC8fN+OUOpb+eu6LG88+EYN
DeDb4Iw3Sx3Xmg/lHgb/X4OieH//55CZx+MPqmkFxcvPUsyn6z3g2Rz7EbRpjv12VIb3XJGTxw6c
GOe6JvA1fC1FagMI54XA/fCem/kchMdoWgsv+nRqLSs+J77M1c62DYkgEouA4/sNfmoA+EjyRtNR
LlY8l91uN6OjkNgNVquR/kJpNldJbbokhMPraayhbElkGrjyDeg/fyutHoMSBYalIrvJIAW/GZZl
gN3s7f005VA1GnjvG3eByq/jrJSck3Wuxlz7DBok4+6MAWKlky6I+I9lp+Dmgv3obDor3dXlX/HL
eBwbZ7cDKWInoop/4nWTNMb0MyzlZn/sP7N3AkSvt/SjyyMVbngsxPGpwMHXARsDmgtYbAJZndBA
jDDpaYc0ih1F6WAb0/AwOyZMcvlsfXrrfeCrlYae/JwANWeTHV1sHB64E38g6NKca4wZGQLAbn5Q
J1s6Fpj91mJdLxtQT+UV149Ks+YYhv1Ie6OX2OitvKbqeDTxQzTAHo9o7Qj3ygnKoOj58+t050Fi
vh7QD0hcJV9G9p4d83gW5xpFK8ybnpBSBaeaoyhUDyJTdssL7pLXyQUxPicBQC7pH/OAFaiVsxF7
QqvDiZoiXUrHLoOyFzWc21VcbNltd6Uc4Y37ZelHPPwEnnl3VjeFKtNoaCukfpz9bUIHU9Q2sM9Y
cbkwfdapjL7DXXxnOHLjLTRlsJu+tysWVqsbxDQ/dRe7IZQdAfXwIXAwDiX7vzdiGU1jLBili3v9
/2axnGwgYsvHTBEn5zPI+ZryQ2ltkvha6a4wKP64KhTDAbrV9ITjS7r6j9Fqhc4RF579OgnogAjh
bXAIr1UMlpZ7s0GlOZod/5DAmR/XwlSjWEdnfeZw5AbwdpxsbcrJfeCUowPBCkGig78VDet6JPav
F+3ByhF/cbMjsUbaHYMLc15uhUlpJyaf/T+Bquy0bCyuEFj8uQT/P+ZlOoaOTapruesS/afFjcPg
CDmAYXkNyvsZ4a7/Nbf7E7PCMylHjCnr9q5nt+6Gj8rs8vc0tu+iXS6Qz2wvpMVQbqA16+aLg06F
q8sbOq04MMPI/nl9PYN/Cb/ekNGLLJU1LeZprqLA44sdvyNkL/xFMXkhEBqMGuPOfFfPF/oPXWbV
xj76MnNItW1X4gdqFBO+VcWMeV9e/jxxE6PZgkBtNVrC8vlItAdSRDccf3Q4ypAZVLyopSgIpaCl
XCTkNCg29M/hVX8OPtH7LlGfK+B2ya3JPal2FWYRkvSpODt4CEPqBN5l3qYP64FggjetuyCaR/eX
u6GpbgPlY8FQrAoHKhQ39zAOW3RI7j2U6vmblEgQ3fXckeJ/GaKa0AtNnvI8+hG0Lh/jXPHIYuEi
pybtvbXEL8R+KhLlLDFfltwKiOpglV4pKR/2qPmqmPBSzncKfXli08PsVvCtpSplRSxRI/wpo5HK
v7rBU0VWjXOqdo5i1xzvP0SwklujzGvI/OZ1sUSnJbYju0UIOzADHD/0kZEwYoKGFs1EPDzEYHwe
fJUqc8YwadgbVT5w8ZJz5cxwIYCrllcR7RSbFmCg146iPRqObzPh4Xkxu+mT4+E3DCazfvwIsAV5
KfRkYzEO7exQqALSG7FxsYnLPS7EvZSPguo89PnnithbI1gpFliHmG01MKBwRp/9ApcWjrsDjl6H
OvrnGIZqejvzNDTylEiEyCHUrojzYCou0LgFohmaWCbZUqSjNiwcqbGySiFyfOShEts+sNpuUVo+
px+SPn8xag1WdARv6n7eOJFbq2+hdgWgbKzL24txgk9kyTKErN/UCh8iS/bZydcu+IDF4KYxFtnC
MScScFQBWR2G8f7Y4q7oCSp6z2zYENROuf8zDP8i4NyYKraYP8j16fR/ZixffCk4yuCKV7fkPQJR
wQO5PaRFau8xhC7Bq9uvrznk+W4ZKCv+SqR6qET6K6cPiP2LzRmvLbBqHcIftBLHX3TpwbSo5I7c
KxX9P4bml4pNOvHCmc7jXXMWNeLFSDcw9WBuK4nLyiapaqp5z7qmLxIEefH0dlYJIvVNLDMGMKxx
4SrzWUj+r+KN78JHi4sZdHiP3/Hiw7GypKX04E2P3pL+KxNKHdtAfVVpdnQJGGbkUIP7Awb1ED3U
x3SjjVXMcIrG/rAVlm2MFEOPP9+waKyb0iDhOTBElultNrliEF47hZT3XIbRBmlfdKoxRVh13Fmc
e5ddkbg5mB0CwrCNTMgoW5fY4S/dW+JeSIyl4TqIHnhdzm89tA5PyKE29/qJMSuSv3P62ppaUXOs
tJ8jcgKcSQljvWU3GY1kbICk6mE+13xeEOX5St68Dug5i8VdWhWhXrw5yee/HK5pGX95YvkiyuVZ
0gK/UbfxOblqMnfglQVTVfju53RTyhCtVoFLSEudJsfW7fF1sgr9G1giYvaTzruVmPacGPzbBlcS
06f/dJJ98Cer5e4X0foyEni40W5Y/SZ9mfOOQC1f51bLTGZoxPcfkgtZ6ER2mwmW/AyFi5XFIdg5
73W0aAp1G2iIDxwSdW53VOhzqiS6NO116RjNxCw8dAIN8JBN4Kll7EArgUOnjP9tYMWzouVkDI2I
w+nMt2UgluzU+7qA1L/heMscl09rjd10nCItKcsFcO8deXIn17ZP/BnbwKhNeQ5y2kN9qej/dv5B
Nz91QWHuAXDoZ9hQDAEH1oTMiKgntFutZvarjpUSrrRmWeMpKpsAxItYmcrdbQhxKgUSEXDdWkc6
kBG5FWLkTzoNf9OYcs/2N29bejuBNtECTNY+mz7jDCsA6JH1xsDk/RiEVRQNgTj5F+LXzi4blZ45
kX/qjzXegL9cWFIdcDshPh3R/2FX6j26fiQICXjkn46+Zr+LGA3yZNn/TgwasE8pMy1TuJ+eNMnx
5VfbblwTJzwjfz8Z8ghvOK//Y+3eCqH7cHxDYoqcqIUexPgKlFhO48Dr6WzVwrekxqrveYX4hipG
HSoIlhWo5xZRYSV2rhCsaOYUVdtzXNJRLJaJ//mr+ZzYkags/o+/tw9wGgKu4EPE+wAU3ziumEmm
btixLygT5oSH+OQZ8GM0vTLN9LnsfkKwdxh+OdW18gT3VrRQatuPjya4vqfW0UpJeoVEA5FACDXB
ilKdYrMPyCZy9RoQYFO+T9/EtphkubE97uPSA/9pd5QWMoLIihQxNB/Ozuh6XdrJYn6oRxNQbeiQ
qmEgrY2sCdZ/LoCg8rejpR+hUVG+FJ+EXD1uoUOTl+d+mAA93oJbEVAwz6DYy8yNvzh5AKm40fJG
Si8g6waE28X+0pWODL8iKeeOhUv6M2ESCwE+WNgYJ0202CV9b7mApy2jXJ6RjOc8O7VnCd8FNSUb
cnMbzFjP76jl74QM1eE8xaAVF8SWJ420+9eVXuMCkcNsF1FQE0KvCKwNF4Aajw2WSTv42s33bOjC
qFaP2sOwpaky5qmwHe8vTl9JY18RuTvHVkQZX1K/H59/Xy06NqaOA9wE/DyqVzq3cYXi4HiEHhlJ
YyOXpemzwloAtv6O4ChkD9prs76LOwrXLboA0TAM0HZL48SMVIXdRq6Up2V5kBECb3Ker2Rak/A+
ceJM4A1psGVxuShZHQ6vgW6IYCjyNwyDaVGGm3AjJ+Y4SpPc04vPra6GhVpr08L2wejU2GlxF9GQ
Fk6OCLBB+gQ55Cu/Jd3U2XmqdmvV9hieoz3qmAbt/5eyGMNCoiId0/ICoe0RU6kr9ovYU0MTSFNU
jNbzF/SBW8XwFZg1aJtmpGuTkVO5aaNYE6Awj/5g0HKfMOr10jcsOjNapUVG1seYDuzmRs3rqCDo
iuZUPdcIy0WEUfkdm/B/VJBwJuyarfn7J8cFxgUK3j7HZA9DF5jVP0HYsLmfDTWvATJAVKLl8pG/
49fQT/+V2dFJxL/LysnWGu/LFTtUAqd9tdCrBqM1gwMY7DOfDAoMnV+7ASPje9tQ5YnxNsGHKCD1
Z8rPuzc6tXfoF2UzYwA7eK+k84bs8nFD57uxjUXF9LJdtcuUtNWN97Q4rsXk8y/tjsgLh81FEElp
6jNGiQVjTHI0FxbaPiPSrcFCWI/c/a3ngojTtPFFI/lBfD4LX62F/JVEQkZVh9DVLfLnKOy4QAw3
5JX6fRc5w3rAIfLj9uci0pkTwRGdmte43KAAocQZY2k4EWhjVRI73zZIVkHxuKqQD5aZ8aydQWd1
7kOWTjRAPVzGAwVQ+D1kFe6LzkKbBBwhPk+fYAy0JN8qHpm139EWLjh/9AmIJPKPMSTUFLqOGv4g
5PXFNeJVtpARgRxYThr5rXWH3mE6lNdPwdrEftNhttkR3koYyvJyxn3H3C6KxN3NJLOpD0NKfasE
YPgSfbw9YtnMJzxDGEZ2HG7aUMEnw3n3j+BhzzGdny+OU0A9WX0Vi/W3wnn6iKrG+okFG4q9HziD
yOEFMLpYXbSAaxOXxvHWUqj2KH11HBGAfdJ96IX/al52MXsAWrXunlHXm5iqt+Dac1NhRBwzPIY4
YeuNfBV0H1w0sEfTleIPw/WgH5uIBoX0m/nBET9KLhSPX+3opCYmczVEG5wDJlTm/fTKXYua0LUc
Hftx1qC8MnBeRFzcr75KBncpz74k1cqFU741Lov2dMlD1EvldoZB9DLiqws09j6oQ9DVSRdhq/27
ffbnNrF5wlK4E+d+nCJR1AZaS2bTjKLg1Rw9pXa+Xeg2wOlLTVMtdsdDHcRoiB86DQCdtOnmbkQv
0a5rq5i/f8+csUCLIaLP7HkSq4xeFwXe479wgyxueiEIBZo/NWmA5KtSLrnswfd3gaj5PQTCcr8G
CHiOgL0PJwfAfwl9dm3g5wo1G4sn+S8bLkzkO9wdsfIDiZ4dyyLqo9tRhSgUZdoqiAZfh96qVtjV
J9ddV6jwxtuIalpsRwJ1LqvDcDbaQ+dZHKS0MG5yzuNkVW2D3rUOTKOfOC5aHotG/+ZYtiN/cNVI
ylzQJHysPJYCfmnVMCjoOa2MHNITuzDyg18VaJdTXuHNuf0/PMpWf/e3uf9Aj1A3mf6M7W5/QU3/
aBMPuiXC3riszSLrioIWBm8IzWILGE+pNhVkyzUuT9ykeHnJCQj4GLlAh71cveggNP9WPSEjvFHE
/izsO/J/9T8ptrnVUjBRT55TQ/mwHGbI+fVHU6scyUl9tIFvC4zGP4MjFPCHRqbULCZRopYXfFog
VPDDf5DbN1zTwJOxfRfx4Bxb3IUr6zaFRIKMg5htCeNDjGWncSWU1hxDUYNWInM1/KQUiMZqq/vl
W24xR/Cn7HMALAuQT6DG6VILx4yajKmR0WDttAHj06bkXktkJKmL9rx6/flFIY0ltTwqGSGcHUAd
5dWvYSBnMQted6YsFT1DbaZpWvnngWcLqY4S/ZtURnuZZ9EsPXeH6FXbb2c+/LFPB85Iqr/5i1Ea
f5WQtTNp8vFHbLaJiP96hGMnqkUlM4Xm25Mr3s39LmFI/y2gDLTTbnEIe/WymUJvzmIwS0bmw90M
Z3CIYpRx2seToxk8vZXKVKmzFRn3BJMAJl0qYtOz/k2jV/p224aCsKedWj//xB9oKj5FXEr/lHvE
FmHzvT1tkfpcNOu3gZIW833qwXQfIg05DVRC/eFoWyk6Uf36pWAnAFaACb5blqfj4LSCOObPvdgF
rgUpsgX8k8Y4MxUR70Vds33Bwd0jTCqa8HS/DmKtheuqPR0DKX2B1jXOlB9Tj2uDk8Cyjk5Cytiy
r4RebCjxdONJamKJp4qiE5vMAoV2cOF66OuBsNbICS02js88CbofHJh6a8VgxSWnOdOzn8nBH2Zb
j58FRWBp1s/pxjaqtWc3RWgf11iOGK3KEgx6toD2J5/eCHygKnF6l4MzWDbku1gp5Knjhnu9vFLL
qCxR5BqiRnJ6xWK69SCBiCCjpsTCqnrOCtZ6M/4kOH+tSHc14SOdaJXsqqAJS7r96b5GEoXdlLv3
lrnUlJQWs8jewH1ID9VbcXKICFv839pwgw2hg1mx4iTwCoMrk/uaz/df+xUB1hwcGqPUMJj/6tyw
DRP73qOWIShCKw6wmF0zcB6Pg9DPl+c592WknqDEp+ASa50Lzh0nWS9HHjMYgNAK1NKZMVSKLz9R
gl1rFsVpxmuE/PxC1NTRhRSPJ6ZVzjHCsJ/h6peRgcqvQrZJ+125z5db9G8ADzpytWRpuutGEWc2
gxuBZsMGyIfdllo8Z8u16Hmc3efseGTejbjt7V56Gs37ldvsGE9vAGb7cfPX7CDDZnQDwNP0mFRz
I5i68pX23IyKWFfSJ8XbDBNkG4D70VeWRwFyNNjKMK8aZwI3N49DsHfHtChI6wTkyKL6RSX2TOiO
nEnq2Hc3QOlsFrQ/FiUwfosyNL2fMpAvxece3WspPgnYyuGvFMJRiAksvcVrOGr9gQeEJ4v0WIvL
Su+p4q0c2DJCTAd5jp8jRyCQZCNRs+4K9XjsvYZVAhd/77gKqkSm+7wqDpUQkQU5makvZFujpDou
xyxQyKjHr1qFxcR6vWATKqtodJUfpHZyfnffw1z+BHvvOmxIi02XMcjwLoWmJRIDPCexgcUCQZpR
B3KTKS/AsMJ7sBsvkWRkm1Ks71tVu+GkT0wp4wJqKXCnOtEHyX/pxkrjVhAb6I4xgQKuuLWfn21P
Wm+HNRC1TyxwzWRvPP1dZvoIkN+h//jQ/9UjEcPGU8mqIAzBGasugpZ/f6kyb9OZbHY95LZ6Pz/p
2wEEZArswJ2K3ryAfQXnrlu+iEa8PRtcwAmuDBb/W2VSjuOe5FIVaVyfkpWsQjLSYLqHxwgbGoM1
1wvUjJa6CJgxMoMDwiN111+ktMd7bEsFMZXylsqtM82vSYoyIu9VF4J0ueAEe1bEeXMqkNkwIyho
PK2d10XpqPGMfvX4N1zjLhdqzzyPcG93Mg19TeCK6YGDq7f5uJZoML36oApohOo0p099uByYEUaW
dvIYlrR66kkH+lOnpNEjDgqkjjWBxQF/yn8WD93lGXakqYwcAto9mglewoOwMhuKAPJUwM7GKyK/
hduzWyRNHW+BP4YT7RkW7kYp3GnxWBPBP4QEY9NZ1UN3LcmzFDs2Ka9XehZrthAraWGInbKkC25v
sgVnxzDizHyFQMK6ogtysWDazxQT8F4y/W+eiwHOGEhef68TNnIiFy2r+D14Au9LdWr5ccFM/zI2
pBTPRNsM2vRFidQy+z5CRnf331fBg0r9IG6twc8hLJxZrUJB6XDNC4Wn68U7I1vV5bCSocAObhw7
9j7d668Tq9a8+CSnBcCf8AvpzBz+/O5xLibpM5CoBM2Bjvlc2uWTgmE+XqXg4s60eeuPvnxw0W+P
12n0iUz38rfiQSgu3NgRBRN74AvWt9yNSEcWVUc3dm7uoGlJs3GZTDYfkwDoV46ppk1820ozft1I
183X5bigfCIV2ort/wrCi9nD057svVPUTZchPzfZrEKtcRx7640CK3t//qGcB9ZIeu/YfyfnQDTS
zsNXMWbpCIF/gC0chYg5X/f1QpC2fs6EYtn6xAOISGn0/abgIGK62H7VD7Riq9wnR1BP/T2gst/Z
BqewL1ip6tSe8mSnYYJi81wCnB98tEbkOh7Od+WBlcc/F1KumoyNwnb21bG/57nFp49O68GBpO+O
cfQWeEBuGCMOvjvuEq5mj/4Hni237ilhozKu2KGViISjURhB8QNEaIlhlW8/qI3XD8SitPRDVnoS
yq2ZCQtr1qJsAcAVCCZ9LjUEpctc5IPJyf/D5pajzuy3iN+lR2GLhl5RTE+4IHW0PlGTxL746g/k
qSO/Blm+PtyvaOmsDFgrZBOcGsCcXkgyZjqHiJMLjHGCp9PhDiEffGzPCI+EGJqqxSsVK4nmLpL6
8xX6VYTkySnZKj9w5yPpblD1YGxfZZJwDrxAthuPR1lJJ5ZbsyLwGW0d3USDKjA2bqHvBl4sTX0x
wZ0RykVf5Bum0skbmfQBSAsgFeuguzIA8mpDiU3AY5Ur8omJATnfmvlu8APzR77HackhoqfxL8LV
BkoMTR8J48u98WjWpxRHvkajzB/wNmcPF2sVet4PLbiBinZstitl0VBXC2yTVmyLVMwJJ2LfRLtw
SDyilBpgK7OyussDk2cKBzYcYMnJ3l5mXAfchcFqB7jGMok4U1hBdJrdGMkwNOGHZCs0wAhDcbDo
3sKtUc6xUgbgX1tGuFRItmNAEt0YuiGNJBhj+5n7h1vhE/QyWEwV51ng/xuYflHZonD2BXflaG9o
ygM8d0Htl+dEvHAVtCtSGzInnOIy+EYuV7dtwkAsMuWB703rk2Tc6U8emVjE1nQOA0+Ist1Z7USu
GiWnPpq8XqXGCowm0VBqex+0AM//9wGXpnqmXeFId7swBgS1zDJlDElXFlWf0yn3oKUNMvgjyEh9
Gm5Kmx6OVwlEiayj7th5UOy70QWC9AopynkuWN39givCWKu4dPh6PpJY1ImQV4W/c0KWF39Ci4NY
A1VSxpTWrEy8zbr75TycZ8RO0vWUJe2SlTYsS/bPaL4MaCovbpFNXz3gtc4xDySIV2/QRp071bOs
ODeQW6Tz6//fmmlGHAq1UkjCIGzwiWydbwgaMW1hv/W7XfOT7LsGi5P5IgCaqItDfdV1lMephq3D
KhoPBjgNwsZaWnK4a11NS0ZENR0FxcwAn24bXHnjl77mnty6L2ExPynVMDk8+XNrU3Yk4nt78QRF
rPC0I1H91oYG/IoJ5wE+JqFCfgpCD8eshnr6V7IuZbfaR8a7KZ4o3IJvBjYKkOmYiS8mZTzhOpf3
2QJGuehXSXycRHPRu6SWHMQlBcbylDwTzfLDZ0IAMS5KLzSTXc+TjtnRnnThE0yNvgnWkhjsg8Ox
g34j65FucU6laZYXNhEggOyGZl9lQM+WacOaNOL5vUtenOiGQANZrt4Y7pHBVWHPSB34qrxKrZfc
0928n6zCGpOQ+LAabwzQXPF80peXClQ+I37UysjByTScSHbWZgWGqEH8KG8NmRVNISITBj5JmWgn
LfzCL1hvweKd0lJLpdSc8aAaXDA/hh+uDBc/Z0ijYZEm60tp9/l3RK1ne6L0vWBgZBT5vvDZ2vV+
GmE/IiO9noMjuzKuwk9OSKvCXurbKUeixQw9Lcx0HNVy7SSvtskGMEJ6o2A91GcxWlciZ6zPdDIl
Vah0iDH6Bgfld+2QavQlTndY6SChFVjWer0EGQHvVeZjWwuCB3Vf64B/bVZyoGRPRr0Km2KqKiUF
4i8GwD0RlbNM1eF2Hz2f470qke7h/AwqW0aMHJfzRTdm1gUN2oGfCV0j6XNoc02indgjikvZGjVK
vmUUcqOQRZ8OVXY/6eDN0ddtXzFE3giXk3A/mCXBELw+9ZbI5iW1ZcqKVmjIi9tZyZYwSc+VKsfY
dNyzFYRMDzPl/n4DRQN/P2+Vsn2bb0Ws+q6jiMItRYMSyHMpc7VWSL3oToB04SnNS9IdwkrYs3a9
uW6yDC21EseF5tilrO9yAU/IWzTPk32q8h/TuJBwTkyYD84C5GEYJumRuoQZb0vzBd7pRAlDXb2w
cIcjLrflScaVro31h7t2QwFplp6qJprjHTex/9oouXV51NxlN+UPwALtIr/kUiCzIGTRkwbv3x00
KHf3Q+PzEhmhuxZWA/7guejrb/1GQ7iU0/CZ5P5rW1/IWGUsXyR+LWBoPU+JMCKIb2qGodDkeLo2
bzRWHU09G6bk+2awDqvPex2K9i9mBt+gn+RZ9Yu/Ry6jduVxFliW68mWxrQ7lODH8DcS2h4ThxFM
2eFPBeyrDuNHr54kFcOgsvnb8n5xORfOYm1T0OzOn7EkrN7G+1QkNFDBsklY1umAWwLsJNwReusW
Sg/1ltVExsnuNJAJ1emR165J5cvviZKCWBYoZ0qAO/StMWETxd5mGITaakUoZjHZp3/hCuX8f2xb
CN1XILaa0Kr2J/00WUdkouiEmb8grAMueytrRscyppTFaMwqvP7WPO1igdQD0iVE8HmG3HUT4Rvy
PMx1EPpkBYP4cE8FWPx4KZEXLENp8JQK3vMbb+/5s+G4LZuSMV2WFeo9flpupxuY1u7Xhbz/Gu/L
yHJJ/1vXcTEqFjzZv7xotRPYg5WlILEGsGu+SidBdhqCxRqiy4HbwBKQvGdnK2kjNplUE/VRiB60
rwEy8gPKDx4Y+4jVLBcwQIfkfhOURxwmW16ro2Jp/9J1vEEEgku13tZTBafXe9ZT/EMRMaxUoXPK
J3ZsnFaRywhs/pcV/LhgIAN/W++G+6HjwRW5s98wL7QsmCndnkGYm/tXbBca+lLmiaHzFYs3e8yr
JE5qokGGLporS88W8tXfIE/Or08kxtMLIrNA2TLnnG/Yc9v6H7fr9PP8BhiessSkVgSjChT+Rqwx
AnIiv4ZpCdU2hwQ1pEZXoBH6h57u3pu7Z90JCdCFp+8ABjx8L5q40pWP1FfFsxi3U0HRtFD1bLRN
3dclXdMv6IZxZ1MKPrmxialn50BSX/rTQ9q9Wngeab4bGd2xiE84zBkZcTymG+cFgz/A36wsFzoF
lTu4o0luJRkQbvIdHojgH035L2kjHAv5AP3bqUz+6w1c79XyaNdJWLvqyAvp7kwGVY1m7dQnAf6M
JwyJZWDbME1+/t+UA6lcZXkv2V2/MgUVAGohZ5C1l94AcDMkAMx3X0TAyCJje9pHfLS/OXkHyIxa
lk3Me6fJU8fCrK5T5Np0JZ9/sNzw2zVlAMJcawfJxCwmDNyJc0Fhrpw9BEUcREVXKwvrWIakkWMi
D3gTV8W865Ephe3rbRcOQcl8/6hopoIqb+9VCYyL8Ax/Hi8e8iyoJqMJO+AsAMMBCYJKvRdL1/p+
OGjtxAvSwIJHnR/gJAkk2YtloBruBLNJNNV/AREpbwDWLLAkBrd7I3JjcqNCt4IKoGv32e60em8F
Cm2Bu2FR6hQtEK+COKedcL7TqE+nl2vO28nNIDj/reA1iLDLAz1b81z9GiustCxYWkIm1xjDxfOt
yJ1XYkD9WHmSB+GfByAmpcOnf2ZMgbCGiQwn/+Z5Z6FAYBnj0xWF8PgMKrPKnhIWciUCMJTU17vV
5zq2CZg2hF0kM72/7VCGE74k4zBn0xbo8lBk1Y07WwlGJs/Vncj06ueuYrndoM9WiC2dcl87gZel
EJwUBc/SA4xU/LdKDdXWaXUKy0dHD9MxHHp+SGn/LHjPOIImfoTMJGf+2gDyHtjJ89ubaaoDuJnm
d4cjhFpGqQNbQ+k3fbPrhoTOeBtIFNlRxdpT6qUUa0EagjeGROCj21/O+bAA0Iw8R2/9AMMDUaD+
EQpajU1VApBNCPfl4pzcZ20oEo07HjpDpqzkcinp8OreYC+B7znfEC/9hzvf78s5QeVd1jYfzkx3
HzRyGk0W0XRv71NFDCPJHWoNS+J2ZCDqWKvOoQ6amVKYOhQihO+/T0bPMH4HeCRZpvOgPbVYbSFs
KMWqdqUtzmUm0NAYitbqh/hr+kyjYhoNZpY485rb/WsZjMCGB1ckqmZhOg7Xg7lN+3KNO9u9ng/H
Ysyj3dSUV89CfNtxcnoCa2LyTSsGWNfr/F0CCTXmucb9v1WFuxgKm2NLDlokfLc6rHLOLAaHokIp
yiYZgedwCsEmT7QN8QkFvsfeS7XAyF9oUa3NwYFG1w0U5FAVIjURDj9etB5qrLj1BkxJnRaJTZse
ywpiL3TIZ3RwDkgT3nTf/GeolT+NXdKCLB5JjqqGgK9UmAjITlnP/k+9n7LPgkJt2bafhI4SZiMM
UjtctKk796UDnFLRqhId0oMy9R7o8OkrYIMCvmRaeldgahLkfnc/5CuvIxpIg8ZZa0VrGRm2MEYD
zFkdXUE3n7gzzfKFtogo6Gi7QlOrEPKzN7V4f/af9WurX5ncEtGWHcbf4rmR+IwTp/J/HEVz00g2
5Y31SwJY8N09lq00oRx8yTS6DtPj47wpLVxtXbwMYNUncFiWaD186BxCTs2PglJikPOEhA0L3JeP
gQTZOjVHvz7Rz9jsyBKZWDsQEkTZCtNbhAY+QZthTesIiH+NnoJu0OA7y6ZOYWja7Ry6x8927T6i
q+CqxTt5tCKAC/+yO/cbVzux1mvO4fnyzrkdgNzWuygdmP7WqRgxENsnTUl6PkChId4A27XpwsXj
f4RLbDP/Nm1ceQKpWrnWA/NN9De60yNmK+l3pTKaCbDxa9nPVOAxUL0Mpsuqh7bsC+KnEv12Bhu9
Cy/sCFqA0mZ/WA6eiuMuNncrTU4gwU9DsLjYqiDY27395Bq4hW0js3g65JXZAFgcYu155mwcfHPl
6F1gVKc5Sm/ACTbF/qmEV5+qAL6Eu0+t0r24POkpzjFu7rg+8TdQQ8QO20xFKrdhbkbU9FmhmkZk
aHaUqp2zBtUrRLQmYtb+J3wWSNIIi5WuSQSW+207B/mwP9pIRx4anX7T0rCZGvZgE2BkcZHpdJHQ
Xyc6vDPzJRDfxa1d/MDmBWhTeg91oAQjdw+peKq4QF0o+7LnpoxEax8W36Hq/uLW1EXzKg+YP2Ni
MgrmnVix1Lj17SEXvif0pVSQbyZps0WM9wcEq7YMyBeChVRhk/+OfLr6CIjSRxlPh0iLOgKUfXR5
yEG/Glmhp8aVNxOMjhkK2PpgqMPKAiKd17r3j3dmKY7T0H2P9+Ns2m/YA/MiEdlz4WXFTqvuOuVc
07SQua3UrEVeVZ+daduforFNRje4r+s50YliZsp2fhEDG0GSCt8METKOHTSb6XdYqzLSGxXymihS
WUUnygUhslPvmDbY72kvqAPVjCOGa/EBb0O4GAkykzwgOA4RyQQPFCdXNIksijAsBj+UZyuEuhjv
2dTYWshapFaEaikzOiXVwK9VH924ruuJmMCjVQPivoz8ORuGOFwbw++6moo4FielVw+v1F9IydWL
YZHxVyXIND81HoPuhAvuBTgIWLK+XSiceZe8UhdaAnXQW0sYNxS3pp0qqhNC5C8/43vHd0alD6sh
8RuyCUo8w30syeixKKL4zQIfDG1COHi94kDwMafA/Add/l7Kl0lw055BZFVbpdfxV4WgQZWmFyIU
qwgYiJ+6pcW2aH7EwOZTb/7aS6WUpuTGqF/HkZ7M8UFvJJu72knv2RDFlFQBrFHRVikK+3Q6g+BT
5TQ83mBOs96Ep3nbWZ5o4xol/korWn0x6cg2AN+u9hEuuofUdGpk7Z63HWpYGaXb9JjU5E54u1VY
VmIyq8Sd5Vk1DUec2us5SZw38AwHZc6uBsm8Qw+bSSlFE0a8MW5oiXBNTxXXTnAAqo9eXalstf0g
bkrF+CsBhjsGjDAn/wMSyp5DCD6Ah/qc4DH3/U+5iRDbf7nB/lpAob0vVmOS40U6Nfn9RVEzCTfO
i57TaeWqMQlXh/BQWJ3bqv0gb6kjOZLsi6hJDDgctu97RD6CvqGoOdBYrfp7/cyEPMBX2teLyGGA
MHuygNHCBo65FKdcqrFb9Hy5CNVaV+J7oniYdQ6ntMXa9B2+VbOF6sc/+x32XR2opnVY03/MpGQD
luAc/XZO1pdpQrLuMPDCK1L1DqafxpNiK5n8cWsTrLdXB8xm43aNkQPmDm8Ow/1WPDC6VsVEw1Cr
4LrN8yqawE+i2qzrEpfAJtZjaNn/+cV976dp1xHcPnqYFlekFCOFgKP82OuTHDXbCBSScTUyMcE9
hPjxtSHFxDY7WRAq0RwIELs8/NdpBV7EsEKLR20IdOjqhtfihoSPFB1IxaOIVX2KqVZhnQGK2Zd5
cFbh5NkCCWg/xU86bv210Bujw0K7UqHN413TzUGBlhPfpBfPyughgQwNRtHyuvWE2CwgcJGCd9RK
kawcs2qPNkasLsPMVC3PyeNaVfXyOfonuVvmU/eHgDHqDfPRgD1JfTr1kaQKuDFpd/IepAj150bg
lNhxt7D5OHqhw634L7NYxh4iUjfvHlzr5L8JRXbrJlpuSKwihx4v9HmBRdZ5jjKvoQALEb/eAt/Y
aIdgAsswSudw6oO9xFZm6B6UI5DWK4imWMfowG3mA+7qrDnY3/uB0XbYc3x5MV69sS0B7D4kXRtJ
ixs8YoD5yOh2znnEKQ7jD3JNzteyapeySlr8icEoC0hJ6p6WmAdZLeJ93WY8axQw9OvDfj08OpQb
htAAtkpKBglHoIAWewBUcvqM5/e5dqngBr6hOJ7kOPCsC0LZb2s7eowrYtvQukrvf0jWBw/sUXDO
MaDG6iw2EDY6zWcwUrkSgqbUPavUvprUx6q7E6VOj0fDJgAKKl26LFZJuG0UL/TtfAa7/gn+NBUp
4sUeWqE4Vdgj050tRk1JEuULpb1W4My+6/Y1W/yWH/+fCcR1yL9nHjwACylOraWAG9M34skzGJjE
xSBKZHLG6A4V861nqKuhyDDtDtM4FocYR2YH9NAPQ1Awpb7Q5vSqu+YiX2On7w4A25BGcJK3URkY
N+YSt9UxqlhXcadHqollLJuzNORRZR7sfbPuI+tVtx2KdSCaLR8iuHRgTldJeiJCZLlTo1odxN/r
TYOIXadBGPh9Q6ZuscWW+ltd1QPZird0HGzSGTSJXxS7epiNPz8kdEcZ+N9l4h78DQnJHq9ME/oo
DiztfH81MEBOJGwQ/m52poHn6ATKAw5Hbaqa4XlOnzcQPGqnkdSsyaVysgz2Gn9EbOus/sY9clmH
U6bgx3lhL/qjAM82KOgeVPV0sXoupW5s4KGOiUxqKcD036OHsPSlD/JxkA7ea/cGjNV6ljYbbV2R
ymafACNE5HylgNvWEaHIwKdm0mK7TusLKRQuxuHE0uUQWzQBU16/fh84M8tuwTlmbYbMJnz+wBpF
peWCTGEllJZhRbt7uzNOsuOWl9IZy8wVGRWh1frKhHcdmgc/qL4bUQgvKLQT712n2WI6fvljVoo9
Mt7ooL7l/n+LNWnCpsLkSiOm9+bPawROY9DaWnuPE26WsRnaniq/S5vhxEbLPU7CToR8x9fJv7tp
d+CV0mzR98NeI5ntDVgRvy3Zu0cVnLp6ERJctMxeJOrgNiMojj+MNUShStcGqk0a7R8OEWYBKmD9
MNUJ9O/g71TncJgOaUvrsJmY2o+u23NswxD2ama4gyMpMsnPg/inRn5iHZq+2HXC9PQ0LdJElgq3
u2wAAXs5yKF5zdfOGOu8uAJbeET8c2fLA7rR+L+cEu4am4N/0JNSMk4/3gNl3EUAwzU7vq6KFb/S
3CJOa6lTf5dqpHatNfgZTglFHG3svxo/XxCkNaBf2c06AYfFPatO01IUQ00cbsZZAvtkS55xMP/G
IKEthg4u239z+UxHpd3mmHbt5tC0mHAj4hTEbOzn5AvDZ4AOCrpWnikZdSB+cqFcMejDJa8jFkWI
3DgW+sv/3IHesNNF8s4wVKd3ScAOv80GY7GMN3wCW7071LCEj6tjZJb3De2F6Rpn2Br5gkOJd7TO
yN//gWxOhixFwR40Qs4fBd782ev8G6w9d0wOJrZkSxWsHsYQ4cvaufxdKXj9Y51OG9F+zPJqIPhC
6rPIWPxO22MHN7MQEusAsknUCIqmjXZCok/LJmehnbFYMO2Nq40HOGW3hV+/H6LQsTE5JIgXUoVc
HL0d5SQahu+gC318jzAOKQIWj1sqgv6eApdVMoveIfJiaqrkYf3Rj4b60GU4gq40gi7niDrOZAgp
XTCpVJvZ1wtuPAUR/5svHQBCoiP/L9Jl8DG0RKM5B2EifIYqffVfZWWzFinW0GHAk4xhY3ZLQJEY
qBve2HvvY3UIWRTL3SXk+8H7E9M+rBzophZZCFlFdvB8kzKO7WFBtb/sDPBJvr5DSAZHhKdnGO8Z
5brtkGVFzpKZSFRGecYvZxiQT2BJ5w5ZVs/AvhnKX5Im7V+9d4diavU46ODvYUYKCzDVzxbhy7ua
pTuT3PSc27rMeY6FmWG0ixxlndS/xNkJZ2ta8DaBq5yJmSQ+uE/dTuD4Ixx/93T/3oyjPtmB1r8V
FdHgSx2HdVVnYG702vxGP4Ht3r1pAqyp1v7/fR3rbZYsa2VuD5Wz9Jw0NmHC9yx9fYKCIEeojdQa
9osdNmvzfWe9CZVsnJOibh4AGfHFvfxeciByGce9tk2R7Gha6CIzzkiMK579cDuRiB/paFl07APw
m9eLnVTStGeujW0VcUIg8/fhUeuvBp2vhxvH+Z54eynYi0oVL1krI2X1xY5N4o34+8oScHj2DawW
gImAhXuNGH2E4FcHf2bNfLln5cxNXEzFz68rMGTPy0FOLAT1PH3VuNqphgIyfvx37J33n9YRGOob
/fflCjajuBRqwrqZwl00oG437dTgbU7SM8w4othdHAc/6MqvikUoOojhb5SgYckHPgc5jfHV6FG/
HCjaRnKxL6I6oeDKZfxTmViD1JtKkRFUsDGx4Ly5d1TZHpOx+H+ZuT0UYaxfR6KpSOUtyQCTevBn
tHKdbYZAYZXEteSxHEI9jzCmK12a2SejvjAYyQrtH0OjOnCs1WqeP4n9YcWL/rcXarHdJn7IYDY0
LARMOqT3AAfMNWsacgQ5F1wwih86wYY07CXHr0m9SJk6tcaKC456fEGXHJ1bKWNx6PcO1oWnUesj
VhYOQHq2vbue8qtVUSK8fzNcecFprGceFnKMslHK7fbYcqFJCqk/fLh/D6OBkgDSUwaU1EcxVPma
ujBpDPl6y3yXGSx12YPfGQNIM1WvtYSBbyqbfMedZWuCo0RNbazUO9vDfQIhQCiJr1F50reiofTJ
8qFdIACAjLxPDr9O2Hv1trW/FfwslVm4rHVW8OIu7/5W9/V/KodiNk4XKneErUNKriajZ6CvCEBK
OL3I3JXUC0u7e340zVUfDR2tjnXEzTRfR5LzaDwfqIgYtYrGmr0AsipmVma9XSG+JsHAeqVLJ700
5nyRCW+UFGhf+LyS7O1A2x6Vz4pggLIVBe2Io4uSRr4kCyNPd2urGjI59g6G+P2kpXvNt11cDfy1
4bLQRprhaHVCLkPQdwdxrRNR9M14kSwgNRQv2ZuRJBEZMui9cgRb4oK2+Q0j/TCOyaolUSxWuwAR
F8aJtMGQqmWq9NAap7aP4iSrmPV/JpiXaqu2h/ah5yH5GTNnL2OeX/Z9qz2I5wSgt9C83P8EvaQk
lDkc8UN2Ib2YJhZOLi3/+UsUTi10xPuT4xwUy9Ynzm0r8nPzct9neYCuMuctReyEq89ZfZFzNI46
FT7G7rod7d9DTc3ugw6VnMUVWCueH2kVUIgsb9lEKyZ/K7aS6ytkuwHkjgsjpoaak1CMWf9frIxo
kzeSkWSdli1H8oal64hQAc+ALRsIcKuWGbMk1D43UQJegK48tMo/Xw6BmZD8p1/UXvNpc/TZCoED
VlqvyZnfxhKYJqj5R5f6e/GTgQ1fWueZQzv5gLBi6hr2pBI7m0r1EyDTyxWFELSZjLz91ULcLPn+
essWss2jVrHhq6vZM5dOl4p7QS+o8mtAfYpOLMWcm73yRbLpbHh2YChQtHLPjeOne2C6uTfpB9A6
7k5w12lnRdAiYfijGuCBhiAtOIs2436VC5+5jJJu3t3h5omiqpzNR72yW0b4LAKTB0igjqktMQcB
n0rgiWwxOsP9X/o8fhhY0UhLWX+oTC/cKippjfHbFuoh2cMoTWZn1xgCeNTIGLndiI3ytNTOGG9j
vG13pHC9/AAwM9/GGq+Uh+riQn14MWcA+ckpk7ITyossTJXFFz+zX9LZOmkKQk1zXwwODlFKV3C1
MDPM34e3X/GjcEF6FLEiHROKs5RabKHzRrCqaZHecV5FsYXhsUhlFtKpAmANsL3cF79ufb/CnOSv
tYwiFm+U9M12x/fPl7XC4a+8ymnbxQomYlznf04fy3MOFqQHpRi1uQDqYVBLp4eH93LAXDsmZib5
eD8E+ymeNi8D0ghOa38DmjoMica42+GhUKxz8UBMFeJGy+zdwhG0WpLKBYZb9JhIydluRm+oj/BI
ZoK58xKrGKmndcf4S5wFiIMsCQ87HD8UY/12oOq+R25dHD+2O7wSxGH07e2pfP/Wno7d+jnU+9HJ
He4mP6yj5pO4CyZO9ZvvsglGOSI9CE4AebU35Dpqo+TTPnAb6mpftyRLVFO0J0OqKgwLe0TPOmzo
miB77MyGxNnvnSMQlb0tOu2fWSJCDwUxo9+F9jVkz2JlFMkqah74Tr/G7xvDcxzD8gAv0CaolW+e
yLB9iRiN5bH/nk34R3/bNR4x0G/uAFQd/C0vhewNd3WNqS3NyCxJIbCP9ZbLT0CXRKV6Ce08ygZ7
bYvdCKrmzFw670vxGHi0sdGJRdpwYrhZ/1/17jtEda5uD5FnLnGQzUb0C8SaAZXXn3jfFZd9ZXYK
Zg/HWVLCAqcdgwDkK3TK7c8dK97ZeRbIn8nYG2B4u5Cl5sKPZdCeegkqcK1Yvw6Kci7rJ17QzOjX
/IzCbenU3dKPxvew8UkR1lRu0+1YM9m1OmQdCxJAjrS2FsZ16qkRWVB4eJmBT0vbJzifsKFw4ayo
m6clQ2+sfztJYwacZOJovRlUPs+pOKwOeh+zse6Ui/60e11gTJv9lUPfDu8sf1NOnGdBcpmDuSRB
tPvZmNjMImpwhKS0T28RDeFtDtdimetjwVuQ8HYcRPfHDdeKmj+QyGCV0S2lZKU0M18B7Bo3tE17
EhIuusjmrkYwBmTUckh2tTrOK1XtpM6mn9Eap/a461JR45nXA3dEg99Xmi+kbAkNs4yr6FR64lpV
3ObEdDKWVwudgHYpSFG8olPV11KGwrhrh0u63U+0AVt+BCLaBJ2ISKa8Xr4zeHm1Crv5VZiYpVzZ
UjXkcPH2WKy0i0kQWi8KGhUc2wrA2lF/7r1qsoHDG0xArPzMKKY295Qzy7rj6rwlq7vt9+1Xcbkf
5pQZy2vkuz3oRj5Hkxfen3G5lCPa6Plmam4w+JyHN+pp06YiUdoJ/L3BjIo3TWiVtrVcxUhH3OSG
zDXfHwo0GHlC4BaqBuVZyxLOF1MnFjGGmbYTogFapxoVfLYaIKdlN6rg9UtP0OweFysC1+Ebk7+4
bHNuUpRU/S0yPc3oxHFyCXaJe3Pv1zNbEP/Vt4fpKkg4OhzD3tEvM7TCZL1ognpncLlCEgO8xVfX
Na/Grw6tL7kUbg23+iXPzPF9xdi4+PCdLj6bXPjrHb4FMXOEne+zZSjm5vQ3CZ2ZZyGxvSHrm8Ci
C1744kCDpx/sCmat8+qFYfdm1/4u28le/Q2/0LKk3lM2amx7aBR6OAh+P8hWmEPljr5tj3NU8vyN
LmxktTa7RlZvHbNcPXIZMbz0aErOdq+dVQ+9siVwcCQEW2Cq6gkNrFMRDVOp+zDMAJlOsYYdGwqT
FCNPyQVf9CH6dBSvOpV/wsDoaHAkGaF7HKYk8XljsDKWLWsh4jLWFwcPjq1kcC7RohwNgwquoWhS
ctdPo4vRiC8LUDEtRloihra1ASK858V5SpVjuZ2xi//PDCtKK7gi33zNnijggewovUsVDMhOZhRa
CKCFc1FUfbTTQEUGzWnIKwA9CZ6V/bjIvB65BpmzovsXkcbXXAveUduqFD8b5Byge2Ntv9etht7h
YgjX2f2QpNSGHiCLcWFCpupMbcAZCpa/ImmjKJ+S1wbsOSjthkX0GX+W7vwYgbwy/nB+8Rhic5T0
2tDH3fvSfUYaIGOCPwcX0MXYmn0Y3YSeR59hxqO4MJ2pvGvmf7JCWBRQtQF/VzPoWb87qxFGM0ut
b9+zAXGooi4yDtUG/VOoFb3/b43+pB4vu9wxHLzKjgqi9RF9RBlrqYz42qqHuOXWjURXFckMukKk
1WiS9Nf2bJy1jsvTbm07w1P0dhDhVv4eu2DbL7x728Xf1KAhTpasA7R+be6WShOCY6+pgtz5I0Mu
LZWfHWQvkZ7q6IzyhCe5NK1ZVS3UlmoN4qIYnaDyIp8n0y1ZJ4106m3idB64YMaTRUtldcaQdH7u
5L1D4iX1ylABi+oY86a51f9HChkVwfa46BsfMXXX9C/Z43rnnB/t9QuxVi3KrqDGPe2nJWhoKX6I
zXus33ExuSJSghyYmQ7DE//HZpsmJ1RblQqBNoFE+qKhKQfQd8+awup3unZDTdIQMb8fFhDYSMyA
wG9HVhiRsFVn9NRcyY2DIf1ggcHGUbokgU1bFdvBMVJpu0X5+QUPyhqhRE655Ud355/rDJ3nzjM8
Rx70I9vEcYcfNaTwusIZKaPD3Fo38gAhH3v7ooQsqXJR+0X89oW2olg6kZ5iqvFDFJN1SUlZV2wc
8aH6OTKTs1VEfIteG4hxZwxUg2JLEVFavApTkFtadTfeR5nUk8X6LksLBgCiKHlKcLAN0a+BlRYj
ROPeTpBgumxU/JRJlr+lZHm9dLXWuhiTwf/spQCQ6WjWlQjX0WTmnRzPDkiIdCakgrdNzRtL9Z6z
3iPnus8yBzjCLpdGFAFIjsovkh36ErIdBFGUFipPNR8f4hkFuh52Ttoa/rrrfjBWfPmrJib22zyR
LX+B6CaRiDXUaAckP4Vhn5bHzk7kodU3cmRBq5+d0ltF9j5Ey9OqKQPZe3ebzgk7yfmsPacJHe/A
LxN3xY1wWJ/pJgxm/G7SbtyM7l2CocJwE3IhpXH9/k4W1OsP+J4Xa7yHAcpEBW+ofjqJOdxqXTzE
PmXqrRQKaCQ2IinyGue0UIDvmXynvaneBJ/YBXQodqTHlUDY51kXP5qzpJUvkC1MiJYIhw97grab
XGvIUyyd+KWBnSmRF6bA9LfdyZ2tRqn8cADMmqtZAzKLNtnF4//qBzNyj9bkH7ANDmHB7ZCIZzjd
d5Sp8uTrsiPtulLGvD9Cm2Y+eQ0dcJu7dNG9Jku3q5bZF75Do16IQy8zbcHxcmZ1i+evRegUGgql
k/TqkweODSNV2xGSrIc7N4LZQs29dpmMITnHd+6V0xxcW/EbA8iFfCVchIm0bc498LB9oZugkgOM
LkUNw20ScZzcGiKzgSwQTxnxcdClJRDRoThpp5gVIH0i/smEmDH1txmBMisEfdcYttZlqEjWTlZF
bcYqJ9R4OQewCAFmqHghTCFXMpeYw89pWE+zQ53RnmH8N3Gsh4yKav729vVFUwkoJyk4vo6bv/yX
xA2CAn9xY0ifoyMchLPUYcsrvcO7xVsYXjTorQXCmfTUMv+0owx9/dcDPaSJOoQhW8EeVDDOriki
P15/lj+xExqss+CrbcOusSp9XGCIID/lbRets23RVPhvp+z8hCYLxr3jQSg9GofahaSCjWzVcOmo
sWoEMhXHER86V38/ncr2V/JfWQmUrXi4F7BGNSONTTX8BjJrnI3/Gr7yMN055HC48JOahONEz5kB
eSfs/i9+Z+R6XCIqocyLrKykVPhe4cobZnvZTzv2d6eCg9Q1+KRx43hppSoO07+MTNQe9jkkobxz
ORMeWyhQdRjai/cxsdMrcjcfocgeB88giMZgFmzUSHn+tXlZRX7Ky2J6BmMRf7qnuGThI52hb7lT
D3qXxJ3dtxNHG7jxVKEpGZU1hubi6etf9WMI22Ve1UMLWtdq/a9uhEXE2cfmBBK06g6eEnFfLQ0k
mDX+Fuc+5mhzLE6WNo7v/RUBXSFW04thYn7ISET+6iGwNSJlsjpikdE2ynv3MHKkG6VEyJiBfm+i
7quDd408AgGEIbkLMgHtx9e7AdGo44K2Pm5At6ljfpWdT4UHuzhAUvpXtfpvFZTvgUwBl+DoGnbG
sqcK1i4tAYgyPYmfOoK3lVjODpctEkOuh0D3AvN9kQK65W91cVcK4/HQjZih4xXsHNXfLHjdMpBP
Dij7tlSQcyWED+AXATmEAYBn2Qiec3LUkATLrQ8TZvlSDIe+RSAKsWYmKn1W5hA+aDnJyxiDpH3W
jY5kk5GCFWXhqNVzknJeGe7Il8fObBGotjEMl8+O43bm6jiXnhrFHFKfrp8ezoJjIIOxLy3WSkfl
fw2Luolrca1aYaoSrFOPCDinT3MmUiMURz0bPBGQkYjARtmbfj5H7WGZuCJjgG+qYE/7EVIy32GQ
UwbNGe3x7xwALCreI9b0krzmKWUu+DOZcktAFxoIMafCie8LWtpzvtIEkCv021yRcQkvqkZW22bq
j08jAjiBul7Z97X9V0uffhkymT9JmMRiXviJ4XeC13YJjghwDaNvMYh3ATI7OSGZ6ZOfAKNOPpgL
svZ1r8R20kdiJlkrCDF0sJ6GfyJhoTYlBHFO7yo7Jo3qqM4GkdmcJmaFPTiZcTrxoBPN4xY9Tdq4
Ml15lsqj1VH3xQdrU0PSpawVR5yCkS1q0q0lTDgTyYdmEnBagI6hEwxvGg6MSrN5ZKXySVgcG6oj
cF3jkZKzR0Wq/8axHd+7oiqPvUUuo2WLAptzZPQOXo9BzldVJIXKMvQZhU8w2i//O7EC0M+Km4MN
NeKv0LckHcEYnEpDvHCc5NH2HAJMn6nwSfF1J4J11mmU1cfaMEYe74oO4s1j/FJsOpNfAbPc5Lti
JmvtvqCDBY54T4/+VnqIrM4Dj6uTMoZGUeyiUtZ+NXd165SZuQ6fDrbbJp84sy9iQlb21UizDMsW
+x64nSgHUgtoRpscxAdkDyBWAVqxAzOUGbbSwSHDz3x31sTAa2aiGmHlGP7zX0lqREgd8vru7XTQ
8gMPRHm3zptP2Xfx5zuPthHtpR7ctY1Nq3S+ke+lVXXDhRSSjh8CS5+fZqOFpL+Ige/1y5WUKx4z
Ta0mHGkjXVvP6C/MHndlREueY7M595uH4hNJNnNEoGzXRfM/VtOzbZ7fHPJCgYIR9w4RTQ81glZR
HPLHJ75XX5mSdGhdmjQdq6mPFRAiteOSh3HNJ8wxQNOfaKnakNgfGRgZxthXnLf8g3oGAlp1LHzO
46FllBfVTVfSHUTtiGvP9lfnLpCTnQCbiaTiJKpOn3H3gnk+eoAa5W7s9PvZjE76op2rRX0HtwoF
vdc+2G2FAg+hTfLar4iX9u0JX4xZp0g/HpDwu7Te6nw3NfyDWhXizU3FFvCpN4poj+Gfm4GNSXD5
XN7ehtE3Dmxe1pwpsrYTw14MbEJBsdkEUowL6R60XP9DevFQaqzCe1erKNv7JyZVYo9CDzZ4yD2N
3HGEgqj1k21VEl0Jt/lNrBbd4vFzHo+FQVAEa4QV0NiGMr0nMT2eWVB2f/ZwmwHcnCULrkbX7FEq
5Ror76nVXOocnoTWx+t3n/3zI88LbgRF8/6czDqNVrC6KN9dkpgYhu1vtUU5I/Vw7ynh/FFRTEk3
28v6BuXnahMOa/DwfHQMf95qG5rVAXiYDzZ20Lwf5t1iX6lEkLGXz+3wW4ldSeBpwvPxHkbMzosF
Q/jTZBLhJ8o2PHslxkmlRV4FAyjGoPdTCL0WLygXZ6oJ6f4WblC6Jcfs7+lT4hM63X42JRK2ttZA
76zr+7Nrhjz9aSqzL5eD/mvnLcRsRRk7qOSjGfy3zOTd3xu58gIjSt3VcDbJhlalMjHZo9J3Gylz
7jJ0q+zxHTUuAH0tEHGqv/vVb9wu5lkiV5IUXVlRxSYw4ZpO1uzTpzYfKT8hCVWdbadS8JdUDQBz
ZORNV6FAbLb/Okmfgx2zXA1cxo3Hw0LYbmj55tNPC3IKxLqNMVFJVUWqQRiKIbcVIaL7n0ZPWCBg
6IOZ690XmxP3Ij81OnpbC67Z03ZJpj4hZwvqaF2QrJJxQxgJXllW6N8Ys/i7aQpM5tHET6+YH52X
rZJIkpi2rIZtXVdMmGW6mg1BkmlQxRt21gHArq64E66FsfRdmqRvX3Lfl7n9Z7vh5Yh2U4NRowNm
bJ7ZC3zbyH66Y0B77A4TR6EyY8wsfRrw0jpO+NSsIIdZzIuITU8O/Z3KmQEo7x8CgYVWVWASg0tW
W+97w2mahpdHqgwtgzKzi5AKVCxsj91EMix6oKUzB6SiETnwhnr3GJoZ0+wYYXcMdDX03jadaI39
Q1loQ43wATH0g3hJUZyJa+EP0IYqs1/42YAuoOXasBGHr98sBXpSp97V9H15T8+6WAqfBmX76/og
uwxEVKN39rdNTGmMk2Aedv9vD2jUNr2nWnx+TL2u6BU4kzYauEZiX/au3ksxxef+4FgM+hbDJ3xF
3ZlVkC1tZ7F6VKFVXZ0zR5pYXz7VQH4fpCaUVq/td+3xHGfYwrNFkjztqtB8owTypQDX5iHkAA+n
xbG97qgSoGmUdPlWSNDpeivrSVP/pUQAooKRPKcrvushX/QUw/57Dg3uijVJ87ZT3ak2/XtfSHvW
AvcbqPh6LJ8FDnnNJeO/8kM3gYBnl3TDc1cYUvNqy7lrS5HVGM5oQOpXPPI5IPz1pqy7RVt8ci/H
O+vVSzadQ+7lKkKEK9IoRIhkUE7PNimbsBKKEdXngKCP0Uf0eCcn038Bd9o9zzZ9biFzioY9ssEZ
lC+4WTA8N1csAyOLcf5f7OXjmG0Y4l+nFL+dbc7k8oyUZQR2jX1lVus1ep4UOyt1f32LqD/Tpq5/
lCN9qjLwlK5MqJ3NF0w23cR2TTALbJYppmRZUurNUG91DL7XKPlv40b4DMG9v4so8POq+AD6RA04
v6fMZftjL7RozylHKnb8r3LFEXNnLIdgp+TrsFjD3QdQTyQqOM5Kkbd4h8a5SEjjXWKEw0r/w2Vh
P1dr3g1RMA36BJyOFO7QehqGvpzmJubVkHMF5CzX1dL5w597kkgbPwId/RbMjF3whO3MiETsD/9A
Vmuc4h/eOjTxQAUGLZ+OrTxDe8506tqNKzh5A+HpP/C46Z8NBOozDycoIJ7yFQO6HsRQGXNibedd
UiUq4yvQfUftlGsMIMkO908DtXHrAQeenJ388rYDxsMFHPmUBUY9qKR9XrXouCt32g5l/qmikHQT
ykOmenidN568VML6+N9hEUOhyY8H9gb6WycrzY+y1O/noZkxTGYWAHDUcp1yyXJvRMBz7Bo/KuEV
84X+xDqTEBtnLrmr9VWAjAA3p25Qx7ftTyUpdnhveOvPPIkkTyzcPbbTv1Wvx2xprcG/YCnmYua3
CRD1Piqdlq9xuv50gTFyRcA3W097uEISuCA+a3Np37/4Q8TZeq+ongCRtHymMLkZr4C+J4ALJAKw
CLiTD5xP0HrY50utRWhR6pLrngh3Va4zGGES0KQ83qlbU9xZgqOTiqK3PbSJJghU63fy1oTRgL/c
VIjNbXl2sk2/B17B6z3OrqvWVCTUpln3ZN5mz8fAhqgLF33RZRao2Hjdc9kH+gl+VYpI3RHoYb2c
IVJ8EHgfQhWDw3TJoOwQBvKIvoMeBtELBYkSrVEf2i7JWwaNA74Ur+OzRR4A7g1OOmp3GBS5C3vB
BBWu+6HrKHTSk1vbB1uHZc43y9XfcFLGfa7krWAwENvSgSSFiqq/iL5tp/a0cpUe9d8rmhGINQly
YmsukJNxVq7zjVHTtERIQqbe2MD3fpP4q2xS3mLweLc5dl7+5+uNM9MERA1VH/Vp1+2l0ibhnyd2
rRscVt3PsGQNTRAlZ1lYfsMwBGAAypyIt72iu4PdkTwjey5bzSTLYe5l/MAQP0PLU1OqxQMXhD8F
NAF6Z/6q+qmW76iwcfUjlaUoQS+8DLUNc6DOvqpL0OU77sOOTrxG050qMY3qX+rXX7nfZsgJJUaw
RqGk4ZlxafeYdRByWSn6zDgzZYqjT17LD7ONQoH0M/TnYq57eEX0xcdy4wreScei/jP6HTpc9s/i
Lea+HBppdfsxIfP0EoFdMn6axQb8le7VUptuM1J6QR2zsMddmzxVNW9zsV5de15L+dnKylJ29VHX
Xu7KXR982sNx3YXaSqdnnXNqtynEQatex6qiH/mhZUCD6L9B34J+rGEIX5hWKoavqn5n0r/Hww9D
huLe102PkOtiGX9aVCGN9TLKjzte6IzirwrL/5D5mQideCzONd5rE6O4QkOc6SGJN5VH5lapRE9e
tNghPpl92c3btOcGBv7dfrmoTzxHug/ELe8E2ASUJXDgNnpg3PIZVZbkg+RppYqjAm6KnT+4Xf2g
q0NIxgjRtWeSp+yHWwT9gZluuClaGfYJoud0ssN+9zrJdxiP2somjEJZY+rzRzebRIvNWxXlNS16
nNsZF5efzpRYswE1FNVq8hc5VuSFShF1o6g0P7vxpKbV1SZvvClqFeq68EulWNSvLmmyv984ZQ0l
3lOHMCzMWoJlNKRR2KGzUIxUxhXpP//Sw1kN6J2yRYLEt5Nm+vVb0I+YxiFULwUmeT9nqOByajA9
4/LjclFrasNTWPJZ6eG/MkI8NIa/639qLu2xMmLxiLIYJ9xobW5XbCMiEwyreXu8MruSOOXdp232
8A7TK0qk813zOuHLiVTIx6dnyVT/gJT6ZTdS5O4xjfa7IhoOu9YjDD+fwvcDFbFSBcrxOrIheXqT
wwj7XXpT8UOK1hukGKutjapBM2+h0v7+yA1vOzYFaYNtD18id0DJ8Ze26y9NAp8/hbiLaBOiTMfI
MZ0/jCEx95ttODKmnnIvv9/f1aUmWJttIG81Mjcn4juCSyR7mjLavEVieyn1qRA2oJ+zl0O5+RP6
tDUneJ1lz5CTXxNW+zQ+Yc7ioc/Iu5fsdFJK0O87MIYFI+QrMrEfDRWKjqFV1/sKq04Ip23aJ/Kz
jftRyKWDOsdveQmj4GzDlOQpCPcoXarfMdPtT7zAUFtVXbURpkHxy6BAbWPHZQ/lNMRN3icuklNa
ms6TreJSffDsRFm8gzKvNzHiIUlVyezb6dIRgVjp6dOB/e+CahqicwGHVEwmjNfSixWO0UarjLCC
g6YMzwM+rBI9F9Nbh1+5z0Ye+7LbvL9L0Nss1O7xN7OVFXBSpIRQ45mnXWe4oRR7CdiS+dNuEjhN
35hHKoQ1OYFNLKqMDZOv1WPeX6sJYvGv2LE9RSHjiM0XVQ0Qxsjsjfd99Yo2bwkiY5m5Tb/iiw0Y
pRM73yqdKo0I/cROZCjwBzHRyyIZp6pmJXR6wnZPfUParib5Mm9XJ4MLmplaoUdtAxo0scrm6zQD
EUsgFx+eu+b3CKgf2NWIH252rB4mzqcfyyNh29idm/oT3tpK/o+Wc2gmXQLyFXokDwij0qQe2IAX
p8RZljjRBhvgdmtFtFY8DG7SSwY1FOkr1hQ8kHiC9Mk8oUQUtOvF/WqYGuQtxxAljEeXMvOMbL0J
aJN+JrkDT7UADvSHARnuDjU8h8Jt4T/YGlIzy5cqb7P3++eimAZb2fGK5vXm1aNVKyfXUe4X4c6y
u11tPeuvo+Qgz3mKIeBNSB2RMPf0KAJ3rcwXyRtoJenYv3PXKPgGdaBMzUN6nEz3OjPvwaZzAtrq
ZFAooWgo9wyKY0hOrjuor9OLgApfJhSyubRD+yWAmV4gzb+M7RWIQp+GWsgXr8sGwLqXFPjdW6G+
0bb/dFM7kh3lkKRAvLg35zgG5/1LLQRObTRw9374+u6mXAZnONxi/N+M+4U2EKDDinEaQwHBoKI9
ZQu21N2NnyWkOs37mJI/9Zc2MX0JghHNu89ukW0FAINgigmagG4DAbGsX9GdJG5Mtv4l+71H9fq5
LRxJAgfH0KbrgeDC9AIap2rZkiK9KChQ0GXpwT53grNFPWY9JhquFqSJXcByshr6vBg7E+b075eo
xLNh9NPiufJwUHMfIb7xLp2NzeLkrgkA/skM5eZkXk0jY1gJbc7bR4GG8gE2AdzgGI+VCBTMrB2k
IzlP6hAFRLkz7ahtH4LptIkFRfap5r+CKRdIw2YhSsQrrhnOxZtnbhLu8cEr5Rxk85F3uSewLDwP
xAMAfgNU3qDj2fbD4B4AzudaJfLO0rPJ1z13I6ZoBGJweMUmU7IsMIY4jA4Un2RhzQ7FL2QUKzur
X6I0rqgsmzs1W9zny1DEZW0I0dRdIM8yTObDQPBgyixeby7EnyN+lUnMtUl8iM2ePPs9voUZzQro
4fZVVheJUe/ktA6DPTu3U3PIrbMqtkP8zYTylJb/lo3Vis37ikvKSihZZei77mbPSPyGyHUhgzXv
emnxx2ZP5qYWdD7Kloc5LkqpOdIvNHuAdelvtWcqC3epeLGGpKrCLpz2lIMIsYPkyMB4Be/wjXT/
5UkvFtB/w4NxtH3QXbvd6M+pRjnhzi7mOqXY+4fWn7amcxszv8ZhI+LO0ZQa9CmehKR07H4IGcru
yQzIJg28RsSuJAR5fiZziV/Bk7quLSNKJnzIhgc8ANZPm9EWsvwOA1IIASL9nEW/c+605TDAP3VP
nfM/WffIC8WNN6EAtAIQpmx8VgsgfNsw8rGO5OuSYCmFlaC8ABNDfErJXhwyEjOd0MVdRUsZMfZC
6DrvOez0SuEqtGvf9drFILByaNXHOKwYdS6r6s3GrLZKqjCGa1cgxTxT8LpgYcYkJUBjNm4dJhqq
kPP3Q5Q1euXyqOFGLyz5ptBGgQrhNfudcugPwZkwc5Omjal5WSUh60qQkl9xn+2SK4FUqNjhcbt4
xIXStrlDQZNIpWeQCwXUpAtLsm0par9P8v7XVeFxMcCJ2tpynb+ts3pnUG0CzWHPgnkKimz135jT
r5uz2FIy3Qax16KZcgwk04VY7R6sQQXcHcPL7yOAcDovkFDBu9zm4tA2wZ39s1b9uXY5t7BhK3k3
v9S6YMpKzDfihcXviQy/u4Ws/aDY0FDndPRX79vYlg2Ts5WTemrsmbwu8+eQfJfTSrvRuTeKB7dj
WTICGDXcE2vNTtA86rOK/zayGyJEp7rbcMft1SlD9zSokiA+PjmlvCcQfnaywrsCslLAc8GyYY30
9phfk29DPR3G4s/jSF8Xg5r0bwQTia4D9R1lPK6+RlLx7QU3XSA1u1pnvJf8ZfhKNEGj8WuY3rpE
NenrLMyKLT+HvdfRHLvGnAgXs37A5rqfJbuUiWNmfDppwnH2vIz/8Sw0Us5bkTvjbXqI6lfBEuwW
nQTgar9bnJjLfdFFvOyEw76e+mCRpDcL7/ctxE1/1OGgLWf7FKZ0C8ULdnrkp0pafQxUtD+CkaXI
sRuAZHIV92M6T27eh3VMuhyJxtc3WlX9l16eEclQQill1TdvNk4f0ilT+mt2eIJ9VQz3mjmIAwzP
+xx2bprKCsRL76NAQ7NYyeykRpi0LVH1TPGyZ4XJx4NvGk6zX4PnOQV1r+5ssAfXTinr1SJYJJWy
6Xs8T7ELToOoQeLlPP7ylopIxVm6Y5WZHTlZL4DiDcv8wwkXVFzXkjn2bvXneS/NIv51DTzWi11o
uu5M0KGPYZvjQnwPJhCgUh0j78WLrelpP19yg6ts8T9xQ97pBn8XMun9tUNM5pGWnObw6no/a/L3
Pg5t27YR1m8Efo804YuIqC9aEDuFgKimVlMEDHjl+pnH9H1BPtv/5ldHhG3knrON7KEp5zxePPVd
zvTMlAPoDKtKpnPKmZXXWQGFHEioEgjQi4hwDrQTr1gF+P+10q3Gm+0ULDOrrJkcBmNSnLDsE8PT
MPtkbqNebiiu6Z83fI9yh07tmSFjF5jnHKeJoNn7umwXGFnVNPViJvpOLUu9xLclV4MLTYDrFXC4
w2tv43qTVy7H3qbts6vjBiC+blSsNaj3zye/3lc+813H28RmJvavleF90CxhqT9H/7vZgjAb055X
sDCy5b4XzXQdC6EW+vsEsSFCz2EPzuAJoLBrD1BPwgVxCtdqoZviKiW7QR+X0FF0WbiHBG/kchpi
mrqdd068c0W8Ha70NRJYmd9azlToXxDHdqRCEKqQ55G6y/fQ/jkasOiEM26knASFytjVgmQpprgD
KFoBQGhbZ/EhR/wN8wUBBKK8nrhLlztnpl7e0/fpE2oA2WwWmG4ADtdeXGXGFC4sPsqF9BVz/xL0
0hXuZwFUVvKBE88djvpRA6LEkt10IXhepIdCU+t6MH0ip80paPmI2m3maGfOrK8askA8CZg2nwFz
tizHGKK82HS2ZxqubE2G5UleteksI/eN9L3R9RtZLhFFHbhnjDy7Q8SyemlaYeLuRhZM8ZrQL8eV
gcSw8eQ4qN8b1EL6+85v/FTmIPkJq6U48bSHgOVAevL6EJSRtsPFUgyUOayKW/RhXUBwT7IbydnM
C6YpFtJ2wKP4GYABNe2od3jPpT/v9FVmAJfENDVTp/F+vAco6TokoeqGE9mOAQLG+ll+bIwdejpt
JFJzxi0xVUN9c99mvViRclB7mthTANYaDWUZGp+YEDY9koBUPuTFdvynJu25RJhdD/Gw/BOCG4Lr
vsqRuoZEcgbN9V3DmhjjVqmel0wQi/8C5qtWrzbsXlU27d5UhcHSky5LhVZyJJA613h/nVoZcD8B
y8gDscQUctaijrrDyhpn0ZSIS61vVLHYtJIUeLhjsGJYB7MG1pBiZyxU9T3nzp8m8ai2tEqzx4C0
EJkn6LaGvHu9hvBlWmOMJfI1tplLGZy0p4NTw25poPNJiIvKPFkgYGdZCDv5B7HXJwpcZ5gAdQw9
r0SnjfHn9Rvh+MXbughZk1n2LFE5nNRcOXDqToNSi+oH7yox3iZQJrDjqlBTYUxz7O1FG5Ok8b+d
OT1LEWrgNly64IFTvU3PuxKhDYldob7vxaVXSOfSclrRuKFHol8i3bzKmHbgtmpJbMmhBXd3H0xU
Sr/hn4NWJ2TQN1I4TeYfvOSoDHXmvxNF6R0Yvqmn6V25STwrw2fY2DeAacjtKnHdofKs9NkzIGZI
jj5Gsb8nJV900r3WQjPsN/5rn1X73uPChfAgSU1tmOPh3e4S0YFZ4tyBfTxSptdl07pE/H2roiBq
o7R99eeFbYFOiPFg2VIoCdbbHLdwVMhVvT4YNw4645EbMlql9DUQLm6m3yACGKamZpthmz9ADcmq
l6ouuxNJjY+xtIrPt4jcf2JELZy/fkQb8nrG685bPr20svz65d8atP+BcxqD71Yw4tb/nBsLL4XX
vrMQA2TT9J1p4qe1DtI0f6ABTLYfBxYutYcKTHR2+uRnGplGkLJz2hDxEqIcAqz0NvcmnRfTPWho
elOs3d3bnd+PM2aBOZFEDVBbz8/J9Gxzol/HSCjXro2nKO4Pi3LogH8fnFe38AoTy4nPk3Ij8Dew
IuH76pyuQ2aJOVWvXwfPffuBafuj5lXbGSPMvOorDweQCRY0ugTXMuOyyLm1ewg6z1+6q43PcY+x
csCmHl81YGTRnjDCTnNyYznAYoIUGuZXg8xRy5KEokee+aopSiAyClLK43IvRlXBAY2NVTXpssQy
4U70cijywlTV5MutEP82cag0OKxnpSFSX5IGauXJUr6jFaHU0Id8Aq6Y2mETaCWWp0c/TsOfqVt6
1Pqd5OHDXzTs7gvPM4lsvH+HbVHoh6Q6xXu24qrm/I3kiLICHx+OXZ0sbx4/tfcOdAabFiVjUDSb
+vuKeIOJ5E8W9BTIiPRbtqCUgIpSApCKaFWgz7crTOToC5KK1OnbSWYSa5Kh4UW8Y/a9MIXLZlwp
hbJDW5f6ICSYwZGe1OOnaJ9LFBeFRQTluQPdUoi37czwvG4ou+QLa+rR+P84I81mqGATDbMU1wvL
FBGbz0m8jKFr2xvlg8NHdO18CYuEqo0a0tE4U/igReYcT7890p8PFs7DFmkEudjUCRtIH/retadT
JXI/Ya9xIEsgaOSeCnnUoKf0E5TAXIdy+2O0H7nAhaWRry3MP9BrzAxiW3uXo44fFls9yureEwDD
tkz3jBYGuag2p4OVW7V/GF+ISGCtQmnp/xE7HbRhuXeQAA08RLoifHZo6yTOYOc97Pn4AqFqM/lg
z4wwJNx5bDgU8+HPx+vzYl2rUdkz/d97Oju6ThrpcQqqY1NMtXpXFJjGWLYNsSZL5IlJIA8hJqv5
7QSlspq+yb16jqgc1Bx57RW0B2STrhF22m+c2/flVFaGhZOV49bglDmr8pwCqZMykkuKcQ1WFsnD
GNKNNTo/gMJJ1g//zcSwSVoIViKYH8PDnwkUJEVhiPd59hgRAol1erSFrB1r1WplnVULfUsgsQtX
pZyAf2y2T3Wp4tzhVdzNYm83LlMytCy8YcysIoyQ5NVonfrj4LWBvnBcF23eLs5SgN8QI/bx3cc9
CIOHHjSjkXi9/nsM6w5gVT6/htgCxaGmg3Amo2CZuHDh5dg9eNHJ1tNmlPy9eh26q0FjqQM7GoMP
UUgeccux0lsMaf/XmOBDy9SydFQae8ddNd2Rvl2fpt9vomE8IdMv/SpRjjPDPJ9QyuFVO9zGTvOm
S8N7Mv/OimiL7Csoe1MR9rjm2fqg1reAp4DoC+R95fRS11w34asioPLq+BH3IYU3MhHl29GUUULw
2MGo3v48gkNeSg8J2i7SkgDMmvAMWAlwRuzqXYZ3eNKc8AYh/FvucE4Dxh7pdEnjJ/RqKg0EKAcI
9pXZKQ+btSlqFLquad+G0nRXpMTgH+nl2v+vdQsh/K/Ay/5iSV+rkXLYQU7x00qGIz2Lbp3qK9Kq
9GL0jSVPpKFBCbRU0s1cCHA8yNyXi5Nj0egEllwUdZMhBXFr7Z3iNA1TbLnp+BG/PK7P3wC8wdpW
R5qTBB4siE8ZwzQ9sN6u9U4mNZnmZAvYVgEwcX4yIyhmDzAB8+023ZjdD/TXE1haW+hnyTwJhQ5/
Ht9++Skmc3Ibbjzm4YyO6cAMk/Jc/4wvZnCgxoo7N1Bn5W3QhviGrYmGa5Sgvkg/P0xxcu4g1QAY
kmcnOGeIPX79EZo3kiBak+aPWQVTVzMhDb4nJPHc6/XAohMW5wi0ACzdBtxFW+FlAbliqRwFTNgf
lpM+UdJx6Ua9cyL2/tniHURWXX0g53vvMVIsbZKhWPpek7ZeniTiI1HECYE5Q0IezxSnDtRf+tv9
wUQMSrVJt0IKMosIq+5UO4VcNWNbrj2pKlAQvaGBw/vW8qileGdoRFwBwgkPLnwCymcIWTc6BUY3
Fjkr0qnkMXzqIp7K2Vn69g+7ShMSAFeQtMJ/7HlnNPnzfRd0BwBdYTafMVlZsm1yPYp3UhmykhZd
XC/iINzbi3zn2LiCY7EzuQu6EnOxqH/0D3/N3L7le2qek0QxDE6RIJqw8cWmDl67WktnKFKO6sCI
Ow6kNqrzOa0/rCjSugcndpj6VhnFK2v7WKq0pb+nXZt2o9mM32LinQ0rpkPrLJG4dfroV63zuxri
MJfE5JuclDrK46Ceqi7qAtCFjZtQf6YIwyoBAXTRj55cfITTevpF4Za09RlZ+E3k1fYuCXDO+bsT
A0MENMNdAuwBkA06E5PrAIdXaVzpPKFAuh+qqnkpJRSs6ork8NQopqtZi6PUc0Fi3tllIbpmt+TI
sLplc3cLrzZP3esU/bpfPRdLqkdp3HgxoeIgl3hcAh393y3W9Sph/DvWW8dyVN8k2F3BWFmxj4qG
pDKOb3mFanvi5DWj/3xnfzXJ/oEosemXDFcUblwYgoxR7urHW2gNo77i/KRtLSCYBL2m7g5MlLsB
7Wf31t8nN1zFK7ON46Gct9JUMWeA0zoDI3F/mvD4xwKfDXsh4UiHWcw6WGY112nDApT55Dat8wsu
L3oRalvOYhk3pFF5lJu0JOuHhA6o3eJvrNqojkUwYVj/U9z1yyGWkI8INJSWsYwxYAKRiXq4qHnq
zoTSMSIxlRAlwvTQYV81NaJJeLFYKYznf4CAUc/RZ+DMYEzFBNNwsIUqZoWCbgaPrExUCuOJL1Qk
X7cKfe9DWRakVbG9o0tov8LJ0TzfUo3WdALM7BYgZLDjHJP7exao5OoiPVQQ8HCCe96+JnL77unU
jn3baY8yFdILLV/rXpNHw93bT5dpp015qSx9VQz+7yPo6IFLYZuk9GVuyc6uckNQFSteEsK4ivtE
j1PsPQaE1mlemyM+B5CWDpnZpiylffaGxapzllqwnOszySlMrB2Z9GQF75Z6Rw9fpCXMcVSTj6a6
r7zQ7NhMStubJ5/ezIjCe4KCicE3peYY+QUjtRTpnYFXtYJnyp9V6ZsrHjJOTuxf2CAkpteomCo4
Z1sCspH9DEIDr5AuVO68OCbcda43hXx4ArM/MiFqT/Yafk/LOoijdqbIWG0XTGQs4yXEnnVqvHjK
GRvv2Z6xk6P8WAS9Zb9TjElpEsx+aeCYPS1561fnw+J3j+MlfPSphewkNyccxdnWH6zooIps7E3m
izztg5ANMlt6wrp0J+CBSCkbrwki+z8c7m/R9AR2IjGeb0OnDaeqEWPWWxrxZffDyrOyvDyaK1Qt
VsgUn0r0ANY2rOM69A0vVX78KEM3pTYLbWfQNfvzJX/6TiSwDBIT5yCmkSw92odV1kFoHQy9s8St
kgTNAE2sUqvPKRzps6peVbNmrbxqqBztbF0WQSQmxae/eHcZQeu9kXFbacM7+TMliKmbswq1aeTh
fMK1rq9jSrehRW1GUNohYfCjlUCJcwLlZEUTgXGsTQdnIfB7EIi8h996e+KgIIuc5pXbpBepBYlC
2WIRU5h1hG8UdJ8EAB0zajc9RiL3z+fRl1GsEYl+gFZqocKVxpzR33PdhTRJCRT5kqu5Orel+g1X
nOaRi8y4XT2/Ddp4EJzzBZ8V9q0ziRNCaSNE1euLdYAbQTYMOApOJG4gvKKWy3nk9XkBdqQgj4OY
k/hmvt5rg/zCOXYLFppTNv8EReRtBgmjyzb6rVwCH2JBk3oac2DL72xcSfWgG8sLOfTfWYC/P63S
1s2hA51/GwMFqDriNDggHnncX12Id99d1RbdyzzPNewL4aODPR76wy77wa2PvrLkYgFDakx4P79v
MOBqt+YLegmq3I88+3yemGOBFx/AxuR/fgkSb5+PpbfVtB/Q1jHITH8Ms5SiRjbn4qTF0Qb/PjlB
QhOjb93f6srmtxf1iY8TKOUoP+vr2Dbvkiyw4pM3gvg8DqOoEsQxhFo8TQ2QcoIChzDsJfOaK+rE
OpNnq2UOWfYO2z9k07ylL/qsOqMgESrBjSEecstmaXg5SaXdDyfeJOew4tz3iydwLVVE03RA8wYw
VaolgFFzzOnpbn9pMEOvmnLI6FPKeoBQ4ELzN5zTtWFHd/OSucICV9kpMM2bt7SqJ5Xu1nM9Ym/8
UmdVi8G3cnAs1v5QVyGhVHJGZwGox9y5SB3dwziTVb0V3WuJqGKNSGbkPFUEE9cdGE3MatqbqXtm
R3277W55SdBRSzQGspcBcQAUF0E3Mm4S/WiPtBFNRtl8/dGdumTD3dWC1ZxxGH3iovBgZmK4iAnG
hrI/VeTNohg/lKTaVg3CuFjKT+bgjgTuIDzzsUzd5fft1p3kxIGTKE6Cr/b5BQz0AJzlHNq//DNn
K5meNMauK1VDn7CTH49Nxc8iZVxUNEjZsxliVZ5jTVD9BcXVOynnPW8yLYqfC64K30cSQMHEigQs
wGf6X4ngvuRiGtLoVD+QsiR82o3PnJWAdNt7hz0TZvjY0iiDHqYpV0uHkZ4piDnk853fXlNV+W4D
FXRjIf8pbjGMWDxaM+Q752q5gRLAAZzeThlw6mJ1IpeV5nIVAMlB4CXuoyz+DJrtre6GRX/VvUNT
RaV1jJNBP+G/ZEtNqHt8lBKYro6rBahQea5PVRSwIYCCtjmg0GPLIhlt/sp2OueR2vhXFtk+Gv5+
IFpK+v8R8xXp2t/dn2ZaWS4+hiAGyl2FLS2qSN6M+s7SJG8ETekSpi+RFY2KURzX6gAmSQqzs3RT
c6Qh63sG7udXAo9WmJ0rzvww/ORBfBKkneSR3W6jeYMILRPwYPhJmrxOUq3cmSSHwsi5juLb7Mrm
rhixCFN8kzBtBZ398MVBu2UQCRPKWZqQm5m0qSTmaf71dyh8E0/ye1X75pLLXHMchI0SwFQ2K2U6
X59KdO8ZKAGG1X9gzQtpNRcfrHNI3ceoV2R15n7d+P5npXWX2uYpkeNi4MHeRkBiUqTfn5B3kY/n
3U6xOzz9qrO2HfBH87/mW7NGXWkyf0+AnOvTEdHGv2jfZ4zEwnT4Coxs2J3aDxgLGvlPD1CFs37z
8xmwXBeGjeyWatGZttuY2UgrVhqVqbg17qNMCGRe6F814b1phtKLXpSg35hjnhYU3O7D8cg5fkxq
UCQBhrH3yUOmQ3b6wxlbw7FDKJaX3YTCWEjP4VPN66hLGLG8R4M+W3tTT9uQ6/ZQ3hJZXRmy2A+H
X5j36t71ITR3owUwgN7Nmwv6gVMSCxjZIuCbT577vJUUrUQWUVAnm7MBkDLyLF6bH97khku3Wium
m061vVcCrofRSXEcBfzdae3HizZJZTwFl4O54XapDyNsmEBFKmFyNchGgrZj4MYlFO4KvqYujLh/
fMdJ2YTlxZgDyqlZ5Ew71pGflxWQT2vKFeuBOgt+CccEyscb8MQlQC8swTWO6DylgsH0Wqr2rHS5
zIbaRbQuVWn+q5ZwJhRUsP4hxhG0gI86HDrazJXHv4eMrYogvbZ4HQza2CnvI9s457PKXbEb2qNX
Q/t2zjcFxtaeSZ6egLx1PByKWcZ/UQkrZ3HFLruji6MWWIUBhPt2FG/74GPZGXfA5ym0s7vkh4YO
o0oLSIMLn2fOX35e77Zy/P+6TXHUAR7aaJ9IlxyEMWCsJIhRVC4/tQ2rJgQ662nQhg5ggAaVm2Ak
/WF9AAnmCgDg0fPhH3t4EJ89aCtu8+0V+x8ux65qSDfKrFohGthc0vlkH6qr+Mhu7s7DS9FjoZ+q
HhQkvhAf40vjpi4WLR31AaHxcLj5zuEA4U3sszaPAJMGB82iPwWsFBgjWSIOPmP1StNmnIpSPneq
YyMsl8dVnX0n5WxA3onuIL9P4bXc2uQhoL5kTISUTdvShNUMdQ4xyeYjNru7dxoSlWrGTRucM1Qc
G2Onj/HDYdwnfFlZN2hwaa3jfNWrd9Ioe6GmB9tZ4Qk8nAh0/SQzCWx6wO+jlN8tDXv2CN/sWv4G
YR/jgfoDMuo7WODxJ1N8MMem8nRbDehN43lx3QxsjTPSKdvMJhFpPfoDr1nMb8UBdZCkQho808Pn
iLs2RMD0Gwtuvwek6TzecmbKeBo2aKbu3dC0iMcacHFsIMzfL5VP6B5oXHDCTbv2Cg+DTuwS+71K
LzMPWoNyWob2MXmpOHKm8P8R4Nd6cj0ivIgLesRGxLeaV4iYMJnPkn0H+eHxRLb+1YuTpKJ8DG5J
0JhIRN49sAsoqoJjLHuSDz4T3IUE2+eNEyLI1XqNrQ0PumFkG2o61jGXMU8gn3iZ26hqhyIQ0Aj5
bvy0zSqESP+VrTS8UIPXm6xynwomxm+EGBspAOq9yKnb9X1sxU45knaIyqBX1AsomYog7GKAyD6m
6CKnsW7QF6vUOLHjUi/pyTZAglBCHqBDcOWruCvSCamT2n5D1fWcYg9CmhfLS4MmBCK9YYY3KNn4
net9aSN2jhp3t3wDnmj5HhjTmsdO8le/UBqYnSeAUDvpVmIDS17g6MjR9gGlfJ7DMk/WIaTn8yTr
awZcxGYI9++iH1I6o3Q6G3MFpvRj2zZbQ4Ic+GSKD9aSBPPVGcxN+ZObqf0N31XCS8PjCnAieQ7s
JaH0ZDvwSBSWxpo2bAtyND5BK5k/aqwvBhwtmdbdBEK3w1Wa7sLHUUci0lF9SCW6AxBG9DDstr7c
HMIZKYKZH8YYxrSQmvImcB+wqF8aQzmDW6Q00p3vKbgDJbl+NCrfZg3vQgoVlhDcMw9xTqN9O8sy
eYVR6Liw4zf7/GC+r71WwzcVirZsNMenOV0PqrGhcL1NhusloCtJCCn+HZI4uzxa8R3u5E3XHBY/
JXlwHCyvDekqSYt6WIBG7YF1GCdo7lx9I62obb5JLcSK0QajZGOrH7JZWJGab1tVMOMnjJnZ52FF
91ho9b3J7fwwGQLP6qNoEXjsAeFsq2Cm5/P59LDvoQgYHD2vF3J+bgGJWF2h+gPrdwl5Omm1GfHH
MWhkrifV1w30BbxIvBmkefcsAD3co+NI0aSyj4TOBlszEUf0o3HCRyXixoh7kCCbQfmosutp8akT
TgiZc0PKYxkMvK8Qakj5krBD+yKe6wFzszm+ZNGpXMmTsz8E7zPESaHeOU8bPeYdjvfyqL7aXEJE
CrXCaRW3isrhppKAhnonP3dhGU1rXCkL2cZA3ecU6bRSHMpUM+pjUoctcIib0dUoN4p0g/FJLRYF
ds2Lae6q985yJYSCn8zPV8t+ThNZHEp+ltHN7BmFJCUTRuU5aVA4MvvZqhs51x5M2NJp2Xe7uow7
OqVE5JDCOcv0PVA4UURDtjxNU4QZ+nBfV2ToD5Z/6C1gZrAagLjOS/E3A8KXp8Kf8SAKAmCQ67fI
6W+NnWM+9lFP+9Twp+FpvARheA24TB2WYzdHsKyv6ShSrJod934EKPyy6g/BYHU6qfn1RqqzLAPJ
qHFo9klgMq3HPSf/TLyjzIHx/AQcG1GWThf1rSMWJEjqVF27aehiuOg0ijT22+bXs4aOhnH86YV0
z2d7cPNLylsAbki7gdlGNnadBfY3c9eG6DVgXGYDkqJIpXhnbh1JtLM8DC61q3Qr7vzkUYVYdbMe
/MAfxk3xHM5iqm7wjPdTekAATsSJ5tdVU2sZSFs1udGFvVartJjeiBxJsEUMqUlQrlRl8yROwjDq
rpfCpuA/TSMycoQeTxGZnSr0T7fw0Qy6nK9+vX+PNAHoNFVDpm0imWXozXuZuGyEtb/KO3OqD4jg
LRM8eVmG5bSSbAPzhNxf07sEvsW7Kf4NKRFtt+g8wQvUx27w8OLvCwre0W4e/ne4SMU6qqNexWHT
nIuLKV+1qVBAwn5An0ceWDc4NoXgQ+sRoQrPc4+BJLTikeF+FHu+EcJ9auCM+fp2yvLYe6pZE8KA
f1iK8v0vKdMkziEkmNRsmt3zNtO6IL6FustiPVNZ2IyRkScqKiXgN9VEVZ6nb0PpHEi9g1bITeFX
n4rO+pJ7z5tIPOgN2oLBHz4Ks9WzbwssvEo3jhc7gLBZS37CjE/SbsFyRuFCUczedT7+hm/4moHI
ooFVsv5lQM6dOFxf5XTySLx4XYETbk33+7t50Uld4odAkAbilY25hmkJTxMmT8ywBKc04P9RHXFQ
NidBYQjmpLQm2/Tc1YiWjMJupictHMxGurDvamkCEt+HbYMHFbbOXtTJd/U//OnPkmz+KbHDzuT8
+Yv3CTNLteiBJXT0qh5QxXP7ZZth68HJqWYKyfKVK922H5MhOjbCKmEGTJL3CWBl0ySpsv0f+pqj
fFuZgx704xmbt7hkOXQEGLo5G0EJx3v/O6q2ljr87A5GTUTcvuUVWjqcj9CR6iYOBMZvjBBWBWRg
GkY6uKwZMoo00hChm0nHlKurdmAc2RjknG7CxzqZIYcgwPAPLhEK405X7WqVvEIIopdUN6hetYts
Fhc2rIUeqPOVOpiFZ0FqBuHJGMddppSn0os5YJs8VuhORzpzjElc/I9qQ3d/moIk+0MAecxL7G0f
BjGWgmckh/GTI13HD6fvK17yGJ5vbfkDemSwbQSTIMzV8dIfv7RL6ST5DQb2TYS/EY6QsQH2MUfE
j0CTaImtfgE0zyh/XUwdkqBisTvOvy9EDbdisSGrEvQJM3l6x+PGb5wx/NtAlW7D6aBJLdpOL1pM
3lzk+b4Vm6odn4IPY77UMuLR4P4RMSdiDibKvmz4ke+Pg0QKRRXO3V4gQygmPnV7e8hbLbJLY6HA
70Z9IHmOU9Ck9gK/S+56tGQiY0DlpQLfaj7J0Fp43LkRaZZg/EEmlFIxx0OdFeJtKsaVN3ASGNvb
wHViD6ecjktb5Ck2PFE38f61TzujuyqAPtTevbOS3ctm5FvNy+9AxVBtlHo8IYVHyovGQXHzWHhm
Q/pFfgc5k1hGPUFkuIuz4aLPl/jTPmRXtutbW+KMvRlxsgz7SfPn5Js88q5TCJG/bVzlH8Rs/EgG
Lqu5ovilUOy0BmVznHl1tstR7VkZa2K29n7tusDmTqjMgwzNyDEV6jxc1yZLl+sHmvaAAvun8xvW
937IhVRjuDQqbVG8VhjrzWThhVPf+9r1rZKERnQs7nqDGkiRX0zHl5+ApUeFrMzAgAgu5C2V5eHz
fuRiAkNWcSC6YmOhifZIHG/vThsYqySL7WahNXI51uvXnfByvHFPHE2zYGUybHjvTwujNr7xRuA8
gVXd5gfb0mfKcVC2CSUj8Annao+cRKSNyBER+bggZdCtk6p+bdMH8yp8juS6tTXMOhkJwQNnkHtG
GpSzlUdx66COpyS8we2+RRgw/+/Fe6daEgwhgiorFYHt7f7OnOmiEvgW2iOYJ1GXjVFO6NTq5uHn
hDxUz9rNTjK8sschY3Oq2tSfoPk9ddkabluBYasDKTJ2I34FgFYeeiRhX7QyVY2vOciYIwWT2ttI
gDt+vLIWBhaKkeYT2aRXpX5hJOBVdJwpOLG8jktdb4bH6I/IaZjmWPlxc9aEsMuYlBTkXTHUPrlF
luTyvmAi/QceNVMyo6LbjuiyIBNmbEDO5z1hGxWpDOfUFUXda9isp9xs/BfTpMdChwLEKVT+/9dj
5G9riANAt1AgW3QdRYCiaaM+zwOFd2eV5l6dApAbFDB3Xt4IsyKtb2lF+RmzAEoO1uZWm7SN82QH
1cms5BPv0M1Yv+tv9GNFObl8Mo1ncjwJu9ePrIrid1UNlvzqzOGZUVr03Xc98sTaHCDXzLSRifxY
gK9XBGHZWJXHeuBCMHQwLDAFlTlsKHJwdYjUtAt8qDW0ZbQaEZ4LuQGO5vi1a9csS53R+1hx5BGv
ti0d8FgFuWWT2VFY424FE629oUz3DiyAOrOmPeNPw7gAgTQVvQScoFmgYgbZm7z2St3qTvX96HjN
1wWsFtNRMPgPT6DFsS2tXoFJh4RLqU/joQ6RsAjOutovnC/Wo69Os62qCLgC5b6oZmB/ATmpGj8l
QrkXekZOIVyV9+WgIYnXj0NfulHrkzDi+j8a1u98pmlUju1DebNgje9kUnRKGHtpNg+7IPCFoPVP
K1VfT/Vhfgo//gWmTsx/uWj0Ifj+7HtVB64x235Jto9WC91U3WU00L62WN5JGfgefarzLTU7IZ0r
6w9+zziefMx7qy2hq9TnzRHOfPHRCJR1+dVk0MCppOJ3nOFyX2AQ8R75r4Cp9A05UXUlVEkH7Y6i
eLCw9m8zzUAqmiM7mndgbMSCbYQ61h3YA1HMX+sIrbZ9A+0fqnyGwincKRkLvzudXv2Dg/4sgsQo
jNamveJ81MNgtD325eNXrpr1f6IamdYk89pIRP8FkL2Jqh2h2zBhLy71oIXlLenjNh/xj15wAZnT
FHt7ExfIRIoyiS/m/5BlBj1l1i+O7ZapY6596W4ZVVS9E+UzMDhbYzjKcLyxny9REvPUVnRV2Inu
QgpNbFppRmtf2ssbkkIipFEEvXbmKx3B/ZqslH5NcsOWprEhCelS1JjNnMh7iVIDLRDfP54jpGr4
2bhQH6yPOqEWdMOvjkavGyKbhmUdzEjmgAJWoryYwJ9w0lGkKHmJ56Xe0vmJ5a2QPOpLkxI2Yytx
kzIOzRS73G6gL2TZ9mgRKYAJhg4Em08fcMfuqydDB+xaqlx92rKOoc+9G+u4+cFYsnl/5IG3IbJA
Irc5SQm3hvXHXoilfStXS4Vy7sihqJowDjPGcilsoEOKd3TmsJul/RYlX9WocGRbmJSSslb+0Rfp
7Flr4/dMO8pONTy1CkBiEtsjtD9xebL9bjqnPThv0l65P3jffKVuHsnx7InRa3lJMvW5LaeyPgIN
UFZ3mx8n4nKbS2hhtf0bsXOTlrCKeCIIV8gRQJJhH3MqeY/i16T+YbPhvqRJhiqNM17PcAnoHoTl
iOtgWG6tsTYR1SBmU34V22b90IhFkPq8UMaTn6wFfluml/ZbHqwsY87dEILkKaVrR78aDvGM00S+
ml+E1rb26vKG3OVMapavs5egMsfbe154XJ/TVs3p9f1jZgMLB17aORsy/OAshCS6M3kkuZnhkONX
ampM/AazzPZX+bhUG9asjpxQAL5SM3EB+4qc1DrhaLyTXcP+lYJ5hcOu7IBIwQEzBPcXwo1hTTjm
k+z0bHFcxKi9yWzsvhVyFVsAxldU4u99cMbvDU5jJ0LuId1cAhrJ5SOQm8vVYyzvOBCwud/vXaDt
YwYSN3BunCmEOoViFAJqN9Jkrjm2zTzQZsJeTikdfk0AfCfVJeJvhEQ95yxtRVNO5k1QngiAVT1h
apby3xlUdCG5nTKIQQhWxnvbsgPIMH0vHbpE+Mi5PjyoH5pEow+u2nk0n8wXOA3ttfOiWtpF663Y
8/yKopJJh7aXjiWZEqPLtPy0G1m6/4XVBDpGGx+6AsV6PqAaahDoa8PJGvn1SCfk6aWVzc7HQzDQ
lBMYz462phO8ipBgccB5FI8CdRiYKBnC96nNjLQe9PhXNqmKBf8tiiADIfNy44ZkUkYzYQhD31Ha
zkgklmffyYNZTVyf5zCbYYuQDr5cMMeHhopb/0R3C7rsB5TNN5GhfYY1vzapLaj2d4gCp3fnEVDF
hmPzA0QZDnrKRuajo4VQJeGhE3xfBBE0PleOT7vBUtimE1xAHHE02lNgkIqFdwXpZe2kXqYaXY5Q
Cg0XdceyUJQXA7S1auR7BYjua89y8o6DyalKnjwZwDOpdBmFUkLy1spksntW5PpR5shUgj7JCrfn
eSqnjhmoHMZHHPoezlsv69kZ5Jig4sWLfLwqAOb98tXpChLMShXgotCZThiHmlaz9CrcWNtCw58j
9NOpKtW/3qzLgqtRVH5XATgVIOE/xakMz9l8qKLX04AYc55keNFjekkoyk63LGgEWcPxNPLPfVZ6
/qJzIKRzE+yhIoVvr3ZZEPyWdK+5u03zyThyK6aqxMYwU3WXdRTvjKHxXpPzkaX+tkh3gx+pogye
SZNedJHk6zrt0RLpOSh4rkjdiAAmgSumupD+i1Y1+Q5TH9WPxigc5W86i/Ip98mwULzkutnpyMOg
Y/tgKnoWwjp9aImPjTuKI/Ch+GWc7Qa3zaEqadRyca4/gGpEsGeJ9CEo3eO4GQK8NIUFrnemCs0m
a2hQM/eVR9b6ALWXe8q1g+H/ZjdXBkQ2I1952MHVDlevJPwGsipX4DzaCKagE6H0pQ2ESsfju8ak
4q6WPwjXjLidR3dYVcmr+uzt9NRiNuMgKN20kI+e19OKlhbsBNxQJDvEpx6bJLhGChf3ulnArSG/
DoLzxi3WJ+Q3qFbVpJdETsyS6KlbjnbkbJhOFsmvMsAyy/peUtO5GOJSPIbm3iT1OSzwPOmefYss
z/8Q2EqOGSnokYqDf16q+eMplZx8Oz2JYIHX+hPYf1qmGisp4ZG7k4xd6PNWdKCIAUUa5W4ApI/e
GokAjvpscoCC0rCMLYqOn6m3G+3oP/G6xAxw0IuloPHAnzMguVOvRLipg56o4hUAS9DaVYptBzdV
tImfemef9B1OeoTjlTR8yj7LzM7AqzIPC16EBhotke8X0s1G9DjA7hQDOmp00izdvEfvSD3b22/a
9x+K2sVXWoPLk2a0FZYMtlVruzsTCmbHlKY5kR2gplmQtIBT8sc9M7zOi27z9uJCHmjk7gpFTCnx
I7zr4fxJEmVakTEXURVt8k57FYQvt69OjrnSkf7yAYivk1y81YdCSWWqdSZABUe3aKaYxCL/rhKx
e5T6DQ9OeeFbVonlqCEff59HY3x6BWa4GIh8vLRfLpr6SgEdEsl7mFVa2yQi9x/x4gn7xYHu3HuA
lYUgvS/I9oBB9D7bHKvyA3ZpkVoWwUmCdBWV0VCoLsBzPDkSsMQo5hHt2KZiWZa2KdaXEWHUz58D
HQJqFJc0y2vNAt/zTfwXry6WU5El/9gifB53iloCVhITeeQTqngEHJ1b4Io1cR093ogamtLaV8yB
lBdxsjxu9+4Oo4L5rp+rbe1d7eiSBKtRBORXjOkihXa/zYkH0E3kUDTvSAX5/YJBoN2JIAE/kUCr
SjNX9cAuSg7TPh2QVy2acSlFvAzjNZuuyhe3EX6UZxmiSF4xcBIOLq0aN5pSDKUxmUMXRMjOjUql
QUiUr7Q0WTeIqdB35rwbg1rLEGKUUjCw/04Wu4B5bjL5EgkLKqHQ6Ae9ONEmi8+x9JiHBPIXNUbc
tQgmY/DtG2MM+MOfVpOT0nw0eW6BSZDBeiAEVLIu/a0+scrjdV+XN+2Ftc4ZXevF090sV0wqYxA7
XXpMjqdLmg3PFXmtDSbcVPdOrozkyZfYHrfcFEt9+wXVKJdXzTxIeRA9JHejJyodxesw7Iujk5ZQ
Y1ALcWER5g7yVrVB4xmMHqbb3h1aCba/DYQYi3A539fODgxEDXYu1+Poo+sVq4zYTk0nupmTSOLt
z2//zkfPDm/dPWi0uS6mAhrY2ou0xBmQdtqThHHdjACv1vBf+tDAaFDbcaZaG1DLQCHHG39yDs0r
pvN4/qNZJCE0xnXpZdIRxG5zh385zPbkdI0+K0Um9kWHh6Wulf7vxAFs2S2T4IzVYadpZHV3UJn4
MO7zHr++4NJ/9ZNWaUqMWlJC3nbqXbNooblifWr7dUhwrltLCSdon32AfpJ9TZTwT+KUanRdkgH/
6C7cKNEKJ1HVg1Vd5M9Jq/eTzCNhQHp1ghqtrJb9SCyqT8w/qMcuerHRWXKm21QXm3247dlVqawv
NYNa3dP0XeOvZhK8qjuKQmUZsJLLyO9uhVvwqNiZLaRoS/pPeQLNWFUooydmHruOky0FNOWouz4S
VImNBTso0iNiAFyQ4CG71idcUkCWRuIMcH1G7Zb9nVAP30pMPhhk3E7yhspI5tZVuhwkmQ5dmdLm
vnPgUr0tGuvuypabsB3bpwNy6wT1zMlKaZsRcdEQD8a1IRhwr5oFlewC5WByg9IDtkF3/yYtObcg
BSBWw1EBlQN9eQR8Bu3HgQI+qKsyhM1VgovCQFQeBz0LfZIfc2FLtvwtM2D5wxtURgbt9DOfK8En
fUSZwYhpz8zZPTcrh9q57PSykej6NIVuiXEGPL04i6leE5ISi8uEc9h3/pswa8GUV4zV7edVcNq6
7ZsDWQ/3QG14cdYrduEaP435GRv6RYITO6VEZNyvLyRuk201DR3fEI7jBfuR+9Fblm0E2R6pFfqm
TyHukJ58H/M+yO9UliZZvXADuQpEeiz1ApaEQUuOKfBt1RBvcUExhWyCGuJn3Ud/mn1Hm57uPhVU
oY74c8FrjCHEwlk+CaHbKp0nNlb//R4yd71sUSfoHWDs8DrF2cpMJYa7KbUQVVFKh47VHYFOk+B7
cItk0iiY1SImHLeAwpmq8QCNiThTziBErcuW+rYotT/EVe1hN1Y1B2fjtuejUfXlynGFFOHIUK3/
lbq2yHCKIOYJ5H61rOlFY9zBw49wMuiyimoDPHikWWjWzmwPAD+ztVgwxUE1O5bHwtppfBGkO3wy
847y5MhKgfJnQeSJY7DgYdtTQ7ZVE/DPOl3WR9fiJjrm/HBsDRz1mwQabmf4owr8HfDMuOL8QsfF
OP0Gf+2bwJbhkUBKAaXRYotmnQCticZOHHPXgTi2BcwHfDQb8KYxG1xFSikesmEBvDFZyeBW/LXy
yyXcHCxQhqoEjlKsjqWOy7ysRQalICae5VgX7M70SsrU0YO3hemwGYqwzqLAcDhBhnYrvcHpBDUU
qVoPkkLbMkVAxwPVGnbVMPfixueoZdM3Fmoi96ZdEO4hTj/s6a07RvtIPm9db/lImLbtiWJVFUnT
7qCdbm1FtTNTKPlY5cqpFpHwRmrLagje3SUox/h5InyrjM236UOIt62onDvCILKilLyVe3Ty1F4u
Q7Rp6wP8ZTDmx9EdcWrVtMM6cdC04ziaZVgttBA9WmxF238lHccc2/tDQVDJkUDN9OGZtMlDgCJG
bJxUnNjwIsUwNxQhgqI/qtQ45WOP52Ugb2ln/Jes9nB4uJVh3Uq8IGtk5vs0gQd0JPA5srZjkfsj
9qphfMd3QBYj/sW04bTVfUsKPamSOvjdVT9n87Z+UAWAOr4PnpBnSt6cG8zLjaIZJYZcOz6VXFOM
MgJf8QXktBCCTIDxVu/E5OxpqqjeNT1k3zlOWHyVwoq3zd3peptCq9pNhxNQDQdu5I/EHFqiqAXa
awPWnkG04ADi+NbSuee1tV4djtpddBN+ytQlntjrGBw83jAJf0ofZP8gYt5JzgksUa0rT5kLgfK3
k71l9GE1NMaRZhMi2XEntRhGGIRrTh/cUfNakBuVpXVsFiWMjuPN7Jz+6rlQ5bWEfYzNYx3ptcql
eBB2ZSvQOwaHbcZQHY/4mAF/jbx78gZvBd1mF97c0k5axIAJbGXI8Dlaj+eGvybEWlLa+HUNEo/s
yv79xummPV1gWJr7JLH8y1js8xGyeaHfKFcjOHmMiALwTWde66J/G5Bq/coPj+A7Kyoz4eSk0+ix
CZxG8JyTN11fud0lNzZQ0ghNbT/hSjHv8X8kYoMvO9XaFzFs9piFOmqRaHlQyClKlbp2nHjr6JUK
HtOZrCk8WnEa27Cizft1ZvDM90+XDTMXHmqlhdFTOGKKb//47hDPmxiPKm3nJnhPEAj9QeSJzNMr
+JgXu4R+6PoamNEdpSk2cYPrz3XIo6yM1EPRKRx8AMoBJgBWNnmoIvpBkzqM9nydeM7TlE2mMqKa
9PQwakJXwwB1iV9N+lGCPzRCFdBepNa+mzoqfHYyyIcYlyjVJqMrf3wGkp3OAIzOhnOY5ycxDAEW
+Vg1+q+9BEX+2vGdPJ7SSERwxkwspxRQoJvz3VJPoNxzlJni5tB57IyTYXWJmb4BG56iyqhoa+gO
xQ0PAeO5Rhp8l+AwNxv1rIGxiV55C/UiMeayFL+DIFU2JOa0z73jeUhV0nJgGDBVBndXStYqA3Cl
hL7CmIcmUNE9vu2yGaTwtOhOWdRmVxtWyqF+/kxNxmxfh9Ps7FOc2An3BZpho/iFQQokX6SqVap5
2TwaN/QWJxfw2ooESWIVOPBCVfEpdZuZ5/zBK5g26DiFWBEV3sLX+mVq+/XLfH+UMAcm1cUlmr3C
S8e4pMCgPYTozd0Y3Bt5tJmzLaLUeHfzXj2yqtcRKKp0TbZBYWYvyBhOvdDYHCPlT9qoMYbjQk50
nps6jCWSkvbFJs8qFVwhZTNayybKSlXStvW2q5fFhOQ4aHfQEbVS93dnGFozEClkDMZ8UWh6MqAb
+1fZHYCK5Ea3hss+ak8LAhFakiIYgXLsC0gzN61OfX6lyr8tLbTERBRZZDSmxIBx+Xsq6i3TnJxl
p9+MenbWH+mvvahaUa18vDtfZ6RW02hZqhqzE6ZdlBTfDY3vVGCQxn+wkzgXJUV0liwmRMM8DfVe
vSrL4qWntIzi+5XQWHYftFVgSwDpy8Wn5kgKE4XUfWMVswAML3n1dT6HTRIx3aAaDf7ZopuCueuU
nJ8dEbEXP/v3OYXpkK81ktGfkM1LSn3yblFhxMjwA5tGt8wZmsR+jp8ScTTx5SQYiVos+oX9P8SF
rBS4zd3cxDlpdDBgJ0TRoPGmmRdr9bYGLhbXXbIDwI9AprlKgkiHQnY/jl8LyWgitUTgSU5b8hCS
HZBA+CcIwOY4XaZ0+0M9JTUhdbyg7OpF5+OnRow3rjH9O+fZPZ5RGAX0XjIlPYVI2IyXrzlszJGu
pJLKt37sQ+XCEHZUz63dT644oW7EwasAs1lrnFnlwVcXr+qSw/5uWrAyYUZmaRgF4d3LwtgOo0Hp
p5QSXAUlZyD/TgRZUZQXK9kdOZXVqlnkVQFP/qftydtta+PooN+LAzPO77rj0Ph3BwfxaOFWAQV4
KMs7vYR4rHj0UYhHzQEwjzeJrYyf3NyWLFqHw22DyN/S7aApzWtxnO7ZcODAI7YELJHXgUrZ2pJ7
h3loPNWvLg20akEAD5Rg8uy8jM/vSYscgucFhEvl1EEapz4Eapqj/fL14qd7QNnpG66KHyhMqlU2
zlWdR6iDVQUw2mxBk2tuCFEN1KIajpfAE2d/VkJwOZ8cQxN9Y9FKYs9HAgbETqu+GZ+WkP6Oozgm
zO5iDkUxAinc0qh+ywEPtXRbi1zHrgguhhu4CN+QzIlchC7SkixlGzhQ9ogVnUrRO/xesdGul+3K
ltzIJ9ZMmdLY1vQOHISkwrw4BuiERU1/3nKnRM5V3+ihOlKZF5v+fvdLKFyMIzebkqypDyurWadf
zufBSxJ1sRKjx+ZJVhbpRvHoIeHbZjodw6erBXnuSMWMjmB41ER/gHbOPbh7U0unw/mupE9MB7jq
B3DqRW2kwNQIQRdqu7l825eNogiIF4IKWtHkhegA0g4J6XceFeJnf2iQu1LiCc4mngssxfTTV51i
LfFVgiJQvDerc0TEGBvfUeDje2JMX7p3kKrkY8RGuOLk7sNDO9kFNqwIBGuCbxuUrJ8h+T8jsAfz
ItHgRm+EtG9Z8Ek8jtFUchR3yXK12awHUP4+DmaFP275mx6yeruXoGK4y5ystHvmd/RhMIkCJ99w
1ccmct5a9NLVKBQ/9fjKCYI05a+/7Xs6kpIuZuRe/uI+cjiPlkEGFSq4B+vhTKwcMq3RSClyMn3U
ZidISQr476Wg9qdboP7QP5PtknPkbDTdiHRGtnVQzezA2I1vcEVqnCv7qteE/ISo5gTWodxDRzZU
uI/Ckt+Dbpw6aGxCECaHp2CqJAkVHsDohkcbiDvXb5YzDRgIz1o5ZEVpRMZnbzDFp4WISpZF21FK
WaUGCdlbE8vd+FHSgoyUSFJ/evVfSdEjXHR3TaPPs8x+CsxqZeNIaC+feOfdG53muisZL0LAvAoj
sMi6ebjkXsRpNYQcJASWfu/e1tYl1hr0FxxECH+M6xwTqnE9wkyWO3qN5wBZTTlw1c3oldwmDMps
fj0BEXLP3ZK89TmKcqi8P6fE5MtouxLrsp5PYcOINr1J6h31ta2sgBVZ5w2t41+MJToIOD/uB2t5
HSOnxvCDSR506Hgoz9J+2xP9Enrubc0Ysj0UCW1XIAFppgKWVBd6xiPKA8xPg+1K8y/cnUdfZ1ew
qP+uqfVwJh1AQQz/3zpK1KR2mwJZh/meRuGtz1HZrhs4+ZX3Zb9ELWZAEIEo6/Vnn7x1LOHDm1Xh
0olhvUGvYKCrgxp2c3px/eX8jWgSldK/ir0EZRDsz85mUWeYfpfVwoZXoZrXJiHjiaHUU66AjNnA
iKFygJYN0xKBQGa8tUA/KR64asQ1ciyS4YS6wsTHi2oToBNPU9lOKxNyEcvfJtdd5+D84CJAYaXj
ryE4iCiD1KUA3o1QXPIT9qnsM+sgCdDyWcon2u9gNNI5Ck0qeYjgGqrMpSDEv/NLx07nu443PBPF
2yjJf+BJb2DsmXPUyYdNbnc8I7GjnoXoodbIVwLfJTAqhHohUwjG7qMuMgpZIDWKuI3M2Gs8w16K
YpE76S81BAh3DIcfW6PcEZSd0BhL2OreAgEffeNbzmpT/aEz4UQkuyxdX7sE8B+mGIyk9uoE5Nq+
lqS+wHPqX/3CwiqHZoUY1hNKZMCgg6IxdOc2SPt3BPCQICNw5e3/YcoSdNZ2qRoMUzchZEhpHqDk
PBz0NAfQeLlVzih40y4isExcpVcLk8m0uf9VDelW1mWrcL/fQGg/WPtAKIzesHICUuHZQQBRLxbe
3Mg/kA2kiHy5s+IL44Dmc97G6m8lgITUsHuICszJWS0OyLffn383d7mI0/iHpl8qfQZUNLvyl3PM
byO09/+kD04xjvPYRgsKXVxyk3LvjUX4cEFBj6iwUomYEEVwl4P8MeDjpwClNRNlll/cIzGts2Wv
Z/LuzIf9gt4EM+xj3QO7JdfeOf0nOlm3EQWU5us4t6knKqSx5dyDIPrlUoL04Jd2RQYcVyZQGPU9
6a+6TVEK3qg9lmXhkHwz5vSb9o9wLkDDOwWjVpSoZ+gAzxLeNhhwGFjGsWbjZRX10+fBEeJ1Fs5n
WwReJIYm+vIk75ILTppg9o3ep4I0g6fEnkZznroxGlZTrmReO0l4vyYP8rlTsKdeay37AfRhlaIL
sMc/YEAyRsiIBO2cURARe9IAv+2alUjY2Rt5QJjNEfRdJ1i6tA1Ph7BGeaU4yGrNLFHWqeRTYj55
Aoo/IwXIWHXW72yHSuq7CZ3bwym1BhijgK7yENRNmyxbXXPMEmAx3WIkd1W3mQ7mGNwyoQmTYAND
zpVxpFj1mkvVRyc+IYANXLdeCEbyzkNzFWGEtJqZIz5d6PWqelw1T5tmu08yIzry09MgnP8od61H
/2cnO0l8c2OyamoALUvQLN/inlmAz0B1S03rDIqHU/I8iksZ/ka24zNC6eKmaX0oxa7KQH6e5Edy
Et62l4/DIXRlGaprCJqEOhZHKysOOY5mGz6qw1o2tsrSM8Y8M9FFkgRVapdH0ELG/GOeOCEBovg+
YW73HjDjKjNDiuP+mNa/YilLEHOC9hEadodE+WB30SwsLkXkDeoGm+z1jSwcndGwRBGV9h58kPqB
cQvNrXJQg4+EAWDQE8TRGS6leMY/CeDm4IAXROQnyDxFiVw4txs8HbRu0a/VpejhDQs25xbHypVh
iba8zt0wZeh5edBHzSg3yDk1k09bKQ0jh29uV2oQnCixHqNUMkBHpWtcxedEz16dGf9b0z3E+BV4
EhsfJCsEHQiFvI3m/CU7DMcwrREe29XM+PweESabZiKdyXH6Puko3p8Xgz6A40qDDd3YDDuswqsN
9+ENeocsGxpx6adxzBgslUyrWZyzhlXfw5sDHiLHnmT5+JA6dPzpt1LFhjpCTg2WmkI5ZQ3BfRVP
rWaNAA62U52GqOubbRNjTQ8qVc3vUTbc8e4FfS2ZwXgz1WCwE/KpsfOgRjZOcOXJF4+kVvssKZqG
ISqtMuqscqNRUD42SVAC/RX8hh8LsN/exvQcYErT+TxHE/dMEtb6pwCHwgHI5CFNXeGKqrRlT+xX
kCChj++yTzlHwxm5iBQpM2eLrTNJwAcWSxLErPv1o0WbwNQpDIWihTk4R2hyab+26rl2IPp6NwRY
Cgd8mU9rJXAwO11QHk/cuWAXX6OLzPInEExNJ6suzdz2n0Tnpm1hxrJNhto66zUc6OMkYdL50muy
U1xQ3A1kNL6Oy3DGal4zw0EOp8Raev/QsIS0icACOKOt0yVOGfvH4c1dAiRSF8KbMtKi7Fs8z0Pj
90gHps/O4z9oIOXoFuowtycm+y2susBqAqUjdvxNUABTfBUL7hWn7GGDjQfqiv189MM37fRgZLLr
eCNfJL2diDyCPzkE+uGlXCcLtBP8sWNEsOOM379lP7Pmjgubmspd7NUv4/5L2R6dodOcGkamsj/2
8GR+hZWS4WEuoJMBg5NvPK7n+uVWJyeTHWD13wijQpWFwX1awD/G8nbjeWazNecgCcpIeLWe1taz
HbiiqiTQNmuvP96NBauWznGr5z81g4EqmUHZoR1QtwyZN9umCdzgYYLDSj6Oh18cZD/OrJlCPUEM
unrFffITQPoTA03F+/DzGAL8RGwGb8riZahTfFpF29+966NiUt66aoaB7UdqdpjBdkDIG5JSfbd/
SZ4SuIvARblaDUdBUDwRyWrCd3yi/Hh4v4aZResErrHbcIawVqa6ZlRWlyyjFQ12oFYQu69Ioaro
dNqo5dniUjqfvlCex3iON6bfiBfu7qPhQ/nbCoWTlKWvAGdAIQC4FO08z2atzbDwm2RSRYMWYZdn
XZospoNPWOvgIdDu9G/CyaY/H8QvAoLytP72zMIPvGCpUKUFWEeTgPNLAGY5dYs2U02AzrE8PSU4
QSU06sNKFqYYHriR1z0vy+yae+h6xNcMw8gy0aQFdGQADYeMe9BZhsXcDGPpSwDz/9yDarFJQvW0
W/teMw+y/E19yatWVINq7W1T2b9+MI804a20ZF1u3E/jSsWfwen0vZ8Z6en9oKmJGbDKBg2RvuvB
iAtOcPkuo2khGo/KLrnvDDoGzFjBT3u+zbb/gUP7N/ZcwCC++GspNCiWOdZQ8YKMWtqJR1z4CrVt
ZGwGZuTeDn6nO9qPKJDucMWUaMEaNmXoWcRPhUT26XN0QdUhVeGZ51HFrAjEXvC5vgn+UBTcc1nB
ogGtzonubGng0ljgGalhKzagSr7BPrWCxHOISTONC+SWEjgfdMlhWn7sWis1hqV8Ad8rW6FoYkVo
U0SKO8SvNmjvDSYH2p4eB3kl+CkFdF//m/7hM5AN23WnV/B9CiO/z4U/Jqjbc3i7D5KUaslT4Xky
Z6eZCPUrSSB8UjkZa8OLQsYbcA8ZfLyo5NSPufmVoeankKruL5bbE/g68VyzG8U+aDsE9Ie6kPzg
QmZYNGW9AdvTOfyBTNOGgR6+FoeJ6DzWUbx83d21N64ZFbmIljUOaiP4cagTJB7NpeOKKseRl5UF
Nncyl0QlLaFhr3GzHhhyfgpPA2VljnHkU9Atu5T8GFIeClBXNLNRVa24/tJpDIQMCXXBYVxbjHnI
PieoInsC1m118w8oreQ5qM1h7KnM/scQPmVPhVQd5wIC/xw08DkIEdviw8pEDXJpVV46F7QhWgYo
9uXtsGFK7yZCErx6zjn4nw/HRemBoOtUB8DiAXOf9RRYxfZVwhnE2IQtHSHHfkU5f42uAaB4DTzq
kMxnUodliZyRmu+sTRQrdoQlROiBBRAcEeNDpsU74Rz7rWnHWDwGzHZEqSTQQU8qSxjnzLdfCKWR
E/n4y9o//s/JGmsmXK2Dtli+zmDIIIHr/kkU/XSa/ex1DyPWWUsPpse3UU+jrzARPd07FwugBRth
gW+WTTCvoXHwXE4yWmfoSYwxSyWwQNQe3PvVyU+cc5zHlW0fOA5mcb1BT9veVwRXjd3+eadQlKzb
lzVeRhFLVhzvgJeRpKN9WULq4f30F1ahT9IQsMIPAQwNDn+vM71y9C9N/otgvXX/vIJsGzj6xdvN
BVhGneeGiuKOg/oUiTWhWapl7xaBEw2PgZgelYoL58YMsiHFefEk9W2m32bEZZSEQuElTYVmsvgk
nZMjI+PXzo2fL/qNx9sbzYnPDP8iVsW2u0zOkqn7TYFM3I89TWjEEp81e0M2U7HPEWmaGAAtTH1J
nCQO4ZJNbnLt++a5XU8FtbkfwwnV71emaGMBbW1waFFAaJp3SjRQIMiYNreMCSKz3EeHTtJNc0cK
Q0c6KTAn47fsiawWGBItlKIDE+4L0ljINTMMIm0Wjq+FJNlNAtKsdh10zl14pgAs8o9MrYQd2drW
keKx+So5u6MtQiF43mn3aT55DKFV2Pwo1ebDW1t8Y3SlmpEmDuYbhuREAaBnFHXfDdXVBs/dReoK
S1rl+/F8coFdwjWAQ85peASuEguqu9f9NN0QueZuH0WmFr0IOINpxWDgpuxfJDPWBCl0BKZICCsN
/o8D4jqGoXt37MHVZG4+qFmhKStTNbpRdWGC6x6Ty07D+nmypjsP73UMrb9HzJLQ5JZ1UahwYM40
E5oVXa05n+pVF8JzNVbEavvOlXqSWV/XUlDtq8KQp3yM5H6WFqZcLQJxC1dpGM8xAQY+Uew4oJwy
1FZ1mYQaQWHx4OJE9Rutflc/REc0A3zkz1Fo50pPaf1xT3OWlk6cBOS4sJ7K6dMjSBcvJ1uJoOYh
fYBovvlsvMhGH77n/iqwOsnzzrAVQC6WHxKaW1UQwoJSEObvgmhPM6xoQSPEMSdvhkORTZl70Ckf
XogPCdmy77B5LDON8yiB2gyzKsBvoDusalAVf1NPZb5B6d5Xr3k1ahqqpUYo6WyWyqz3zIZExubl
ajMJobCQYYb3MSN1tpWzbPJTLoHWch6bWZGzE6F1T1HWDmT6xdd+FDUJyu9w0Fsi5yggrZwaAJkP
uRNhkyL1QRtsSyD16V3iF7M2ZGhs1v0GLnDSMfS/IZiK3kuEwsMlPeRWtTDNWORPnXqrVKqWMqks
lfcWhOcAEIO6K3PrUQUvcWHM3Ojo56F3fUDZYVD8WHaY0PeYnJZNJEnmmGH8f9Q09/HbiwmX493D
kW9H9Br7giYBZ/ANF3kJw1bJPsbM66KzbFd0l9efXq7Gdo58AkVSGD1bQtsraFWCrY8aJTFnw6uz
wuhXhHZav6/UwL2ANyca3fIt7bN6XCBDZGBkub4wTN1wiGmsGUVQeOXYVRrp+dlYhKadEdrBaSHR
tYBhkHYaLma1q4fqGInDcIagqBQnt//Ht8UNo59OuEFMAo7Mdr0xwlpSnXXKctChY9UnqPcmEb0d
B2CRVcOBzd9PSoR3XKTMWVgfGG99rwlpVRkonTWSrKGOBAC8uge8zVXZ7x7Z+oeHuXsYpU8YC9y4
/Zpcuebwyk1jGYL+qhksE2XtzIcQrSFG31qcXwt9CSq03sGjED/nK8100Zez8S0ayMCd1DqIPdPJ
fs0+gRv8oHCWf3Smdo7gLytYunXBXuPIIosiS5AdMGOMlhc4v2shuvv3IMIHRtD2KMwFR1wXN/iD
YOxqKuknPkPQg0lytjKMWkdNi/RNH+nGlNNj3Fw61UmmGbKdPh0CgVsTxD8Qx7VJ59KXPZFKGHyy
sG5yD7VQyM8e6YzxWFL8AmAcX3JYGg1hQSQGiB44hsH1oxka1ctIAW6jTzVdrBbkfeu5kXF+NHBr
6pZ6fZ98k41QH8Oj5NQ9W49VJknPShdbkcb+nwyOogOkdGKN1cHZDhKkhJCIgqJ+19myNvjx0S+5
e6zW4POkBL9i/YkFIWvT5vAAmH/T5n6axIqlcJ/ADIIkbUDop/6mtPNu1je/zGzAv2z5NP83WS7O
mz7RPTIJ90K2E4X1vRBWsA1ERWtJaeJBV5gNe8b5ARtYEqHCY/AIQ87Q1YA6Pu5O2l1HwDRQ21Yv
f6HEE2XWDqqX/oD4H/KUwp3xZ+ZeU+2hl5RqAYFdj7/DXNvy5Nfw6rbacc9MCIiR5tX5thbBXt9E
0iAJNLZXSvSKbuOiOBwxE63KumfyvDOm3cHtLDHeYz2gK/DD89clO2opGDyumc7a/XbREvsSX5Gw
fudDBaJN9uf0+Fib0JMe51y6tK3sqy7R8TG1LI58fpwtIspMgOf0jzVGEr5isc5XVV29PXxBwNBk
Zm+ftV7WTttv0gXaesUbtEkDkB3m0gMuGpPcgsLL9NRwwedo+f5PpE3xatyO4BXVY+c3ALOk/0eT
KVaZyU96p9V8MgCUg4sIiHWI9ErE3xHF7CL2o8+7jrtc7rbJk4Dd6fvv2DVd6XJooWXBcy/Ccce3
paHMdMpkDIiE6bFiUeBWyFIXNzuKLjukTgS5r0bcvps5GVK7P7XgkmDmn7aIqpJsZLlJx9PDzG5A
RTCASYE9KIZuSqEG4n2/Y3Kjs+QMYC6RSrqdATJFQezacnrW+HnL+sZItpaRNIi5xPYvXk3F3j0R
fMgV+UJP24V11pBF43DHM+3YhYiDTIBVBUP6r3M/cZ2qHinqMEHESMPUAZBqWSbA/Z4C+owLf7Cl
VGkznUugChjXxmKgMaZNC+cHFT7Sxqqahzvhj/KS657Q5Hb7ByCZ03iNuKFB0JZet/dkoTeZ4UCs
YgC2EY+Qal1L+QTd6INiQjmmtWkMG7OKxU4jZCKDmUI1Mcb24557lGKqnAUkitwI06MWUtChUJQv
z0D8YVQo4RUMcT4hNLyTGcBUmJgaFUtnP+dHHBbIAmeIlW8wQi7q1IZJD3r7l3F8CYN8eCy9bIZ4
4rqqwizdhXIV64VapP2Um87x6PSuKbapak6uIUxPfHQFHD2OL2DdH6JYKM+FlC8LXMUid8KBrAi6
pk9/4mnV60WbY8lk2U1n8A/mm0QaB0TyYcNKtflzytMTNPFNJljbLQ46br/cCwtkJbL9PqUpH/hl
VnlqFEi99L+EzB5kEJkBMaC6YkZ2fforRTjKl4apDBcxdKuZnvLaNM5r/PbgmaDRAkf7+7XH5AVI
3FX2odxltnj8cl/YYufV6nJv/MNV3ZWeQnoY1OJGT63PBk4tGQKn6q8ppd+NK4jLn5CPwsn/epNI
rkXTpV1KVdqkd7wW1pPhkBev4rBxU7TDVeRIZ36D6g7Xhp+DfybCbSiNMkRM/Ayk8XtPoofqXTkn
a8yN7zUOHxWnXy5G51ou+E+vrp4D52fQYQgz3BLr6FsHAAq9Eb+X66I44NVMCcj8JeX6nNUc/dQw
PX1DKqSMaAoaRYrbzC9WK8uF9KKlW/lWl2dcUTs8Inc3Vg7ca2DiL/D+WKP0vtmqw4It0ahVM3eb
wOa2Yn78ypRzkqeu7cL+i93sBbXbgkf53XZEEo8DJz5SLOIcYmJh00ysY44TlT4zQgmatyP8h4Wj
fVzZisbroR4fUnUcklYqx3mKus/FK2covHaa5GF/g+OTAxop0XN2Kg4/+Jj+zBDuKzvNTANI11NO
GUntb/+zGwA/X5fQDg0xa7poU51cqau0lSFyzaTzHOmelPix5QStTzykdaIbBGWzYiH0MIR5XwTI
72ZzwqwF4+lWr9pGFA/zVgjfdufMDgSKMSE2piBSZdYJthnqfbUxOcYR1rrEvrhREJmLfWjZZlDK
TXEJsHGI2P99T7Ggjs+8Es/1jkocK7rFicbUJWvyxZKCdtSyhyVHSeo8RZXbneleLnC6ekON6S94
PFd17JERYOogA4TDj3/ZpQP7Mwm1Im5HfgV8AdL1+m9uVeUDhcz1w6fg1C4SpCWMWcEHJ6OXK/j6
lr/z5FBKrcGf86K8S80RhUyZ7WyACLQKMFcGTU3DtuMpbVpsxloCG/a3oclh5tSVibajB8KQ1a7b
ZEZGQw+oKvhvcpHJlc891sWmULRP670JhKRenRrQYbFjT2mtnFiwhQNnh7dP35Yr0yGDpLzYoMhB
xpI9K2NTBzwBWKCGjF1tztdNw8UgDm4OgaZwhnPz7b7GDFA3A5DkAaPA4chPelS/SXEhPU/Lz+j2
k0y5J5U3RJrf2RWhiJUj7LD4oM5b2vS04h8/MweJMyu40mJ79jfZe7hbD7T/kr9zWtUxiYcNhCcN
F9bZla8s+p5JrI3pNOmTFh9tibYGSmoiB9nEYkk9ojbNVMSUI+QDpGGO2m7dw34a1ev/rMVOJ+u+
7ZfCLNxyhVfyvrOG8QAIwneNpIfseIXtu/jKJug4YyHc5WcicCgiMBI1QIkfVnc26BOInpirTxT4
pvrOJyxGMR8bfNSPPTVUjBoyobuBt5S8kh1Rzb/hVzKz9NX6yR6lBCLy2a+2jDoZgLpw7Lyr1qcS
OJ+pX+AGMhiK40/NCgN40PV+7O7DFoTk2RtQ643TOW2iEL7ccsZJfn+9c/7WycicsNRfZaTB/daW
u93bh3gVNCnHRYnvuvSirYEV946FNRAp/hSy+VVflUML+zJA/34MpXsHSlefk3TglEOuC3qgF1C7
1tt0ayM7Ae1MjPqH29Fs5C5YpmmYBMlCmbpfm5uJnXSyTI94X0fVpuI10g06P6ZKK+BI9IEKBrOZ
VMthUocKZ1EDg/bXrC71ce5moHkGkY050GLNOVHpn55sdr3x/0vVkL6X1ns+TcLb441x49vPSoGs
U391p8sJV9PKlASD0UgmEd7CMjGjMBLppIsp9f4d77aGtv0xCfXe9Piaf7Kv//HoRfP7kYKh/xjH
rUuEGPbp7pZyazdk2P7exbsrSRfkXpV9tdba3ZIfGs5oGgJakvBcaBwQrWDKM1Qhsvz5Wy3NJFz4
XAMZaFJGL2XFZcqcBfPH73btwKkRzpw+ig1w3prYbKOepvaj02i460Dz6nYMuj4xgw1k5q9fnPGV
56ua2yZVEPaRMryWpu2SB27UnooJzVmLbPoEG109PUQdr7skRX+lrc2sLoKhrTFrDzjiyUplzLIK
HdoPbCUPIWtRVO5lff33/IRLM4sAuyLkJO1OmXLV+zVv6SKnfzoOkmFK4I1Mw/oNe324C17knmk4
dcKKFF9sO0WWt2yISq3O1z4/GIIqNfeiYqaSJm1wtJU4BTMkWyjkzTEekoy/FLI1edWRSIAkNPdR
6KRFp3Xz3s2JDOvQWSyAEyu17s4t6swZlTalZDRYwnj183hmk8KqiykGtk9cg9qHXFgs3r21scLf
CSKfI+XMzUXoqulqvRD+9JE84py4W/TC+Q8980gMZVl3iGh3QSRn819Sm3XJ0JEpAkqhS7H6lx0A
XQbtZiDAjw2rS2mkJj6EUmj1xlzEjFZV52GGEWmsg9mXx8FuzBBuUn4yP01OrMzG0oSJCdKCN1SA
qYmWXtWUksp+6wjfYBmQQ26X5Y+iawklwiMBXnDj1/Pf0jq3HFwktkP+1P4sMt2/i2c3mm+ODDuN
DqQvaxhbt+dgadTF3NQd4HrzeMC6F7g8dQccEwCLhQyFele5P7wRI/IsmlO2fmaJ8HWB3Vi8lC1U
bRZutIBE2U94YQFa3sLEDSd/7rrwFJA7PSOv4gwyLSG5h5HEPPcjORUsibLnWEOzfh0pao8TGqxA
k/BclGEb45T3B9mtgvDtx7Ep80SK5Nn8KM57ct0HmUwaHFVGfOR9021wamueOs1avlPvaSFSqtWk
eZthx90/a39NWmGG7mbACDjdqG+GgsjYMZ854uLHhCx6/KaerCW6DQvniVqp5HE5R2oLUXbNoS9Z
nI/yu4+DEYfrDCFglYgx/Kpa7NtN1mv6fmoqBELGsa2Ol3iEUF/FNn2Xc3yHNFSStaCY8rKVr95S
pE/49UJqJZaySm82fScx6tPUhyGmhnqOwQ3wY4ETVUEjwOlzzS/s1qms6jtmoXk6ev0WERyNbGnY
dDHdtxm/GuGQOKYuRtllGECTQxWvsjhYgu5QBrvwNXRzQdh2fvyUmVzvjtXKaAJiqoxn7CIJCnMv
Gc2CQiWkVia/lgp/r8lal+aUI5WwLTJ0+FhCaCqJfzro4n7oVV5WQtQ1i5g9sHqUQJQZyplsEgFF
nVjgfioHSQkyiUy6hVhOYclsbHjNHKaK544IZ3LjLnsqmjPIA107CKp60YB8uyoL/sptNQzuJFms
Bd2ApcH/QNjmHPA7XN86fX98q9dV0IHNjFjjQdFq6oNx9kqNFDbBhXdqj4W9LdsW36+cAc9mRA04
k4JAfA3S1+vzXa55BlVcVuHQoJyGi18rVAfF8YK9R3t5LroUdjW/gZ/Dq3QwWdjaPlt9I0pNwDKL
qWQELBsKDjPBLIbsLMrL5JARgA2rcEPqQjZwPONvPuQWv26aMYvZ+tHCLAsA+5QOiAZ+ryoqmzeg
f7QvS6/odq8gD6sDuez7+SrYR96UXHG76sMpZpunnibeWXQjNEK9f1Hs/jA7fGyzROe6O0OQFmAZ
B6PnVHOXv0TiSaK/XHk95hBZbRMgFZWuPfouZjwySvcC3IUYd3Z4WfKrqoe8ito9WyM72dh+RPm3
j5XEaZMJNuYk4ubZBrLUn2r11nAsypvD70kyo9DbrRSSp/m1XcgTapJVl7OFdcri/T/MfRcGcTWh
+nJxF0BOKcxm+/ZzzbWmA2/w1Sa6VsTX9bW5NklIJgQVWgpPK1PGI9vsvhuiXW3gANKslU0vKxe5
XQKKZw8VAnDgtl8kZV+RU9ChVNoRpKc9RmN7rviMa+YIIdrAdHIh5+ZZBufmOKKCEKpGeiH2bUSW
Mp55UMW60dzekM95ATPLhoxsEIQL2uhmIhu/HVxTlkqaKwfzjgLays3xlh1hAiKSh8drElmE7XYT
5Bjfn9GIFrDFwMXRSLH/ndgkd/APN4qiMmQnCwZdZx7SQ7jSavK9XWsAzD0ix8q0VaJtEvCxiZDj
3VSX5yxTCIQjYHEbTmcGkmhtaiYeblCFr8acdb/h5G/cLh/pKmTpzV/cQII86rF4ASVU6bzfe+KK
ZPPiMBRfn22dIPknC3K8f/uyJd468u9Ti/gnLlsaXGJak76Zr2slJYXoJqyJ69CwmIXL5lwZiK1h
fvc8uERBaz7+VIsXROJYosveg903s6Ob00mea1zPDWE1J5QrExHqrbzYuKdDNK56b0HZGBBTXSzI
b7XN6bzzf4hWpjuiYDa6HG9RRtirp5aC+8zZ2TSS2v8j/0ZrmRVcdIR+J3hOiB5nbyG9sKErg8xW
pRmzBdk9hhc7kxbAElSAK3hlsJhB2Meis0rmCVwbKOnlmpxEhKs6SOSPASPl0jJTfn7K3EbjzvG/
jdUESqILEqpTmW20XzS2ZBO89i98hl4GCr8jZvzWx2AS0S1o9hePwXM8OHcZeFm5uJ474orXr0w6
TIha3lFTMcyxQtPAc+Maq4izioCMaJxTRgYkb96NjoykpJDwcvCMWp/iC3gvm7v0/va9I/KxgmUm
91m1TYqZK/KZ6vOkDsSA7GYNz5hwXYxp1CUrsCoUAsMAyxx2nCoU5hegNVOVxjD/O5v0tEwhunL5
ZV2+8Tyu9mofzkC06Y7xC2V/AfjwZY43xwBIbMYaC0F8QfXEDsjF9nY8NW71PlEKP5/c7WvMDJxh
NI1yilN1slGnzHoHdumcInhexT1GWoNaxjWe3uDisFBZ2h3h0sqgANBFyuIeCGbCQRR6Xl38Xmgy
tLWBGIYF6GQpxVx6FGuz/jrd4e1WkVpDWCBsOthuRw16eCBTUtEG+FhCTZD6y0S4WmjGsh4YGCtT
KdQ9p7wbeIyh2siQOH4nc4fW4ZHdJJ0SsDJKXGZ3/mDhwiH+kFJPoBq1OYVbe8Q8UwTwhhrKN/Dz
XJzflUZ4gFG5eR8Uqn9oUb+ZZs84phUYRRyJpbdrsYEjY3g8oOdMuH/Ov9/FMXm1RJrxFJqeqh/i
rKbhGDApGkY8v2DSk6S9Anl5Udk5YIDqKv/amUTF6CXSb8wlN8bvFx+TGLSgONCQl/ObIqk0uTNs
QN1w559hxmu9uZYxpX2yc+lE3CRokh4Bm4ez6+ZQ2pCI5QwOPfQcl9jaoEgn0Ezdxx8Af7oUtxlC
pldUF7Mwh6iPkxVrREixUCHb9AAsXnIPRBISVAJv46BBCwTbZKmdZ/lzEZjbrsXmU9BehKaD/5BP
iYVUJ7tE6AvnMGhQ5QjyndobPDaSGm0M33/p0qz3+a4+v7C7f8NErgRwp713AdAPdCTNzXJUGj36
CbqhJAyPtLXbE4WoG+70jSEk3OVYWl2BqiCd2k4XWRIGoWexI42YisaH+3JbKpUgvcrsFb+C8ueh
nePp9LU18eWD6GIFDYk0QFyK4ombfG/aRDPTNVohwLPEEzTYFpbe+Du7bSTeW+j1++0xHU1wcrIJ
yqioNtb4YjZsXmW+errSiRlCpnNQENaEFezEooqpBhlIlFXJAJu38D+jThDq0pGbuGZHaMZlfuer
OsFGNjOJpltJ2qiutINJMSqYLYLIISAKBaBE3ta26/oOjIXgU3ap2IHKmpV/3LiJ8tArGntSxCt1
bb5sotl5Apcy5PoeQJ6JnKQDbFL1Qv3lLMF/pPnsEcHiUDOJNtWB9w9687FtKQHLiqskVc099GVF
J8hH0l4esVUAUuAaql5h0alqlsqWYCasEvimFzIMnhFiR8wdvHxkQ97ItOvy3eefDLfcVYiTJRsN
fRFRu7Tcbd12jQEH8lC0/EEBsBwODvuPIJjKa2rHiN9fKQrcbhFdUNo2tMAi6+2JSJbL51m1KaB/
NBe2+BFuBO98nBNcSUSy65vX05yZ7TSzNPmDd435LphuxteUVUXRAzCx04idUDSbBhnJoh8KajHc
4yeKDNVvs+1b7m0mDjpPap2OwC/ykhpegsYpvWbfY2x1m+TgYLSp5uarx7vh8gfJSh/c0ifWelyF
1MmJK8dnoHN7VqanUsZqjlR0AZFEfSMQk+2+n5h2ZQ+qYBbpKc89EdsSsOEQRb7gAk9zAFFQbOka
4CnOpc6izSI9tDc9kwXRkVyYbKIf9IrLOCTbobsdQ1+HHe4k8yuLocc/koQzh0swbYQhLQZQLiUP
LMtKOf6SNDNyYs3EYr3hY6QQ503+EaPlSKhLSk4JSWUEKE+IYBPcdyj3tdV7Aa5PLpwN66AQugv3
el65BIR++DbUV4wi9Eott/RAwCE8y1ateYjWgZnc3c9buHFZRGDov5vTFFMoBjErRG+cvb5mfQsC
Ymz1m4Nn3AdiQVIk9q9/FNz+U5QKV4uDWhkGsLIlygCJtkS4FUVJrwBV0uItSZScXVaVjv5I73uB
khwHibwqHyaqLb8kQRmVt3NJ0Ifi/nXcmHOpYNMwdiOWpU7c1cUYyiAl9ytarPuMK7ULcqgNv0Pp
ogFTgwFw5dZS+n/ySoq4/V0GnmiiMekCXVnN7lme1u4UjlOv+df8jukvDXTBcQDfFkN3wR+x7dzu
BdfrKmhgWiyiujlLaFO6mdPKJMEYT8AcGicJRAnWLarmaTmlOyxDKoHhIgoRrJHJ6D+LSUTcNTNH
uCHk67D4NuPeB9A807CSRbdaucEZswnzv7ST03cu5TYKjw7NWf1MFA40NaWONEwCRsVirSynByJ5
KhpwRpc18Aj1Qv1vxvI2UiCseuGn1i2IR+MgiB7rvWy5nroVh0qhMkG7wgqHzJHwcH6LFw3H4qDs
mmi258rWnSAi1uVE/pQzwWDc+6aDVHM2Fk7xbGGN3lngtlziljb2o9vD5Vbs5Ygf1YXXLAWYabBI
QeGS3E9SaUG/gccNYUWd0OJDDS/2XpUbfSQzAuQ2uhDpFa7zRQ2cpvdAWC9X0aiY+3w2m4QhbyI9
1XNNn2qsXm9rTGV4gFx4BBuSTphxpb1Ygo1eZJbhzGFEujXAquPvj+2dzluLUI5aWu+IO2dT/uBy
RwNFmaKcV5mC9IsXnhzHu1GThxyU3zHT2BGXhas9ma9jYRiZyOgZKWFsA+t0QHoaB3BUP8eyajWn
Uc2yaD7PFL7C80xQpiH2qIuBqAxMKb8GLAiD/gKuIfErP55idxRJVZ+4Q9LA0QdBmEzvgQh5qdmb
ZHjD3e2WQp4hEp6nhNsg0S7NKogodoMC61lR1rPSojmtuUgmwOaZ4BAH+7d6qmnbCOX8/WGu/CAE
StdF+LtZ5Wy90vBun1U1btyL5QY8FhF4Abfj0DdEnbajPm/zl9MncbmQmncdJBHTYSL/VX7LuKmz
KyscwAu5v3ivZIl/mopvimOZRySwmfvzrWj1pIfVIlWFvGvrqKczAHuzhTSONZRBRcioH52XaTby
P5LbfwRi+Rv/9a/mo2PDt76NdzZo25TIdZiJ+6pAERY/Ux6OP99MI6/NCFHVUNpTw/IZam23hMmO
gOVvWkiIzrwZRwxPhZNnrOr5cMEUbIckNXHBRUWb6P4Erd8Tdf02hGmHqowhfkqa14GP92ebkDZO
ekm+jmzRrkdPEHk9Cx2EtY1QUUynxxeqEeE0UVn9fmnFHjJEohfaQhAMgZV46Gfr5kc1LXrd2Gu2
smM0ibl8zga6mXy950SH3MDPilRivF3zO+Q99vqvK+DKYX6UxDbMR9LamvHmwmUwagnGvi1cJEKM
Ti4VtBB6lUJ0Agvs5m0ggVZ0niRiupIIC0DsWIT/43lmx/hhPuPt/Md7lAZt4uYdbC9neA54aLbp
Vw17Mqhc20r5D541wTOLzXGT2pVXW4B9rhtQhIEBVxnfSycr9LJwbGGf99LIatU1LSmci8IQx/zq
UZlONLPe937hE/6r14OYD5LOpfcWaY3wf/J9bIQq/ZnK3OL5yboVdwB2HRc5JtLMMjGQvSjBH33b
sb0dPtThIrwNjJSgRURw1jvzHVa/ZxtcdqfC7Ng0RFB1h4WDi+Fg1FEAAaYDfuyLpHBhWbVqfAt4
7//NnzOUspJSYYkyDja6aQpBMRHsWUSddeUq1kDTKH26qbVmv0Tzet06l5l5U8FgxuyhqK1/0Tw+
FN02mWNFEWHkhquuMTcA0GWf224DGcjWWa7cMZ4UjwyMtYqSmhdf0BnSUA7dyL2xkqAc7/CyU0oR
/iqMA/4fUnGqeACD07DpylKIg5mUXyyI1UvtJiqmWpRT9igsFxZv6zScQj4nxFmUk41WUzfj0DM9
67k2/obNQdjD089EjpBQlKr5FMXdv67Zfe29VeoMb+7YTtdXcefTSjkB7P66jiZfCoTrnPd6JVxQ
GZmQ/8QYEeCu11h8BK5MI4ABZuMiAFP0dszwjD00OjdDxkQIC+VWKNl/Z39jKVXkZrYTnLp0+3If
K/143X8YAFFh0Pjt6iGfQo8pJ7ozhSnMiBpWD7Eyq3qIs8TUOO8wTSan9VjEW3IbTDrwyG0YzanH
hzjfPyG+WlymILF1XF7pmFSp/M10gbJJTP7xgyzMxpjaDyIeNeMluVVbd2XcdlXaDXe4FrE4scZU
F1nuJqcDcYO4zieJH/oJFJExCCUYHwC5HdZsi2IpWbiJtqFZ/EBCOtH2K1Yfz1Dk4aAZkJO6Dgq+
RAxY5nVow2lbp2vO7y7sNTe4120UtYvFnIxDHxR1b0o/GCG6ZN4w77vx1UnIIBYiNkFduu9QejRL
JbpWolI9KlyceEv/Lv21sjRFmMXWj257qT8cVqP3ttC0RFagtpe2hyzTkzvZykEPL9WL2kq2npzn
BS5SrX/4G0fxoi9YPIV2sJiEcY/KqxT0BeICV9v14N8T4YoDwHeDVlHsB3p2lc7PfWjC0T+sKRNh
wqBSD7GqcG4pKrPnhFVPob5gzwrlZ1kau7kkcXMG61ah1kTP1lMpWaPsLUvGx7rs7JDeHLqxmMZV
KNpE9b9uBsuzYn4pugxo5gNpKz7KN2Wo+TUqVpZdpLHKLd32dGf9CfAQE3DEcakjp9jB6xTsjhsY
5rWWEiXUETHDSnwcYc8b4UJLfJfDQKXZ3p3i8Wf6rPK154ORiQLJ8OfuE4WXAAOwouy/gbnPOoH7
fDemXJ3uM0JptXJ0kdEaLVTlshhkiHRehx7a9iZBqHQvGeUsNxkjWBsxgVQ4LHo3D8+pN9uM74tS
/g74ryRrZHEw/ODOxZMLPMUUy4csELaLyxpPBeZvYoSL/iHCow2rvt9GEMASnsrG2pLglqsicb2Y
FGUskMXH1UTVLucG7iRupgh2owRy9L548BeQbkw6r7MRcaMGAoltyPzk8f5u2LPK8f3Y4339EYYo
/9tVT22dRt9R4ptx2tvvn3Ec14fOkPf52XT6D6+dcpWjEkkEqv0hCzmqfQerExO2JP66LaqeW26S
Am4SRTnxC6CaTAtOUX5K1gFKV7eRVzia7263AytQqnk5mWowkJ2wanrLHDvtjh0zxp94G5egh0Fu
pJroHxwGsPcz7eNq8oKB3Iq33xN70RzEPHhssu6TbiIwBGp4XoviuY0mGcc2RazCjjzCHnesJYRg
WcvP/ER9KnuGkVy3pXEfeewEXjnsmVr/TI41R/79ae1wbi5Q6yfU2PsYZDL2ShRFJfRLhnbG0wRn
iU2Qm/Vt7Oiv8NR64DyFdLoroZtidt5jHNa9g7mOUchj5nFKgVlacCNTSg21Lxjddii3/12GJvi3
gXhrOd/KbuQt9YkaQa+uS9e2DSKHxHgLSx7ZJ9nO3Hof2lDZPkFw20Scxaqglk7i6MGnqo3Cuws0
rIfP31odvxmN6NHoUBkX6vL/fH/g56MdhDZldbLi8MzoUd78cpCwg3WaG3BhiuCUaFyPByHPMIHa
ZTULvq4UMEgRtsAlzikgJ69aSxpEETqQjTIMpe9Fhdfqq7ftmZkHzz13/ilNQdB7r8ZS7AltOwAu
OO0TfaGC1mGrI5KCZh+ObW31t/RdoaiEwsL4qBJnmya/RUL1oj4v7VoCHIN5qx5+MA2Ix6cBIT9i
W4Zakpv8SKEUl/rWi6WQoNJWmVwiTV6CPpW/tFGefwpai4ISVOzJyFbIdTtK0ZmlzhP2j6hvJday
KqVMb6FNNLU2eTTH6pNQ79yA+zV6820WeqyLzZtEfJfmy9/seLRCKSPKGgVkTjy/DDGE+sjr97hS
1I3e7zq9NMJfgBBI2m+r1Va2/0YWi9CHWVSxkfAqBsR61yWvCdGZxi/BxHlo4XBr7IfnI28dSJCC
2pBrt2QoeuSm/H+k+m01pzjCgJzdcPxX3zWNBFgxQfCF+ZcCbFUIAEnw1kdJHr6GFT6qkEkcV3rO
6tqQS4zxVDH0X1mwnsvRGJJLjCcYrRC/7uGzORgT73g8TiG56h8EPPwDeIPdgvOJhytXrIgdho3z
OYEOQcxLb3+Zhj7S8S0yrE1r8kBWCYUkXUZqFSelyywcG9zlazFSSjlcrZLoCvH1tzo38JZXnHi/
25Ft9PD11MKNks0ggz5QNABTUR2SlXx+7tCNPrzqAi3h8nPCfAq621MIz6flJUdxCYWoGNUNDP94
JJ1eWgQcWB/fZwMODs8cByBGNr9moBNnaBnA7AInQlojsP1rFsCTx5+rJ3MVNkvfgqVdnJFE6oB8
53z+pJJBqLR47HrE16XJ6/WULo39SVljOxjXaizzhQfI2ILlIdBcrufz5L0Tz04VYkmeFX477Mp+
wCaO8Rzkhkt12Z9gpigMH+ijYRQmRisT5E0G+dWIFpE8vC7F+WfLZDtWeYOfEE1n07ZxCL3iNl/r
NfFvCttfHiqEVoDmakwscYnGpjHAwVq/KECJIvVnK3SCUeggbS4ZqS3vUWnH/Ka/ntSuSCwUF34k
erwum0S9kUwOqZBKUqIVlOB4BRfXQboDyGuFRNT/MrS4Tu55Lse6mK/qua2NQeUAWSPr57CrjnGv
SN6pw581NoHR5rM38OexyHJ4Ew//tfPKF16arxTyPRRPkOVzYt3P7QzLgtN4SRQsvwGKQBqyjKU/
4HpuDPq9+G8FfLiL5zZn2UbXv535ObdWJ7EGux8ibSu7Tqpf6ZR4uiV391tr8dNybHVWf3wd7hia
kod+V67Ikm8DQJu2PD/EgCkHry9OawVhxC3YHzrafcOeHCZYd/gU5ukBBMd1KyvZiEZiRrUY+klv
eRTErtyL/AiJk5y0ASy3qpiB9HGCGfk/CDDGScQ/wSWK8r5I74Ux5Zv70Gmicr/mMyC3y2AMazcy
5Ij+E1EmHtx09g6t8hhVIuTJdgvD5fJrCAhHQnTb8+Zcz7l8PedLmyEyXDTYd9wzAYMQMHHRO1Uh
sf6+em3MjQEseptIoMiMak4p4NytOw7vYLCGtKHMEGahA1+J2jD2s356O0eLcvWho3W0kncpMyjs
zZqG5iuC0P7qNsAo7pOqlpFWea4KK9BIbhLK857T5AD5habqhAXhm167IrKQBfJOWqgoYwUPqFze
6SWOuk6/AesIcTdlpfZR5vGjqNslEpffX4rzw/tV22QQA/JMJ0or5XOBFm4N8y3p+JZ2RGa62QSC
+xi5+7J9Kv92JNo4XgZN0G9Dw/CDwoa0m+lnQkUAGiPUvs2ubluCkL9+7b4TyxB7pexTeyZy0xq0
5f58Q7Gondp0mcgBJgLsl1ptq5GfDWggIKoWzCHgxo/PkcDfJrpHXl5O0oPER7wiq+BbTBtTolDh
Vw9pkZE1ZaBPHBXLRZw/UvAs6k9k9WLXA1o4kZEv78SYH2+s+oBaLXIqm4AZ5EOL49hH2bxi14JZ
7V3ZNOZrMhy8DtZIDK4LV6xAom7mx2BtrZakfydoaqPDMUM3xqor6b1hkiPBkSyMDpqGpcN0OfZk
3BW+V+/ezN8ffeBtJuV2+ct3xkFKK4bh7ssRIGt36cohTEiAWDbFDWt6pADEelOqF4O1xfrCzX80
9/vGHy/ea8O/ZNsFEF8tmfymkTTNC1KU1AkmVHvE1mSUQlm2qtMmPZSKPye74DhmMxycw4ZjScVW
F1NeE42bEi6y0llOm2YvH2yKpwdrsyWxegTEqBy/lxikU0v8GLVl0thlcDJeHveEybU/L0wktYuJ
FfZrtU7QE+CoufPZ0M2qm9MP+YniIuxQNABL+bBVUt4wNEXW7aJiYpOfz0Tcaq36V3u/DRkXcxXj
q+ytps/O8Zf0lk3Mk+qEJzaBsx2656sNqyCRKafkKRo5DIiLohHoWsTbtdOwCwB91S5PXTh6fQi8
kYrAVhkdAjKusX19kxwKky/riqc7zrZYQCBy8MJ5vg3gnK0gSktozMP8GXhheXnz5FI9B4MTsT1e
zgmPl8algNJczMwhdTj/kE6OKIxFPoDzaiN8EP//8/t0Rl5P+MAs9g9emiM2t8O/5xUaaKw6CHF5
QM3RXNgvGA/UzMEZwLAYxcbQm8FV5fn9Tk+0Ybz09K6W/P+jb6rTvW4ITsCKwFkaZRbfKUnZMiAX
esO1gqgjwH40AJU2pYwMQazmAp4n9c/1vtY+z10/qy8fSucmQLfE7tOsRIrpLCDUuGEGPMgVQGR9
dH1g6RGLYg+DxhSX83G/qecU99yGaf+0HP1iZ4U66neIejuJnRk5+Ucku9xA758N+MuOTVSNxAL3
FYnWhgQy75etAzhIOr6zO2xLgGPYckTw04f6JM7RmY0DhA2lziAiFPxSgtF7k2Y6jnCW4VzpOPzN
xb8Eo+0nYB1okEGyCnR9ZoI5FkH2g7mYsA6cEp79TAVRfNQok2vh3hDsD7olUEqZV59JElznKgIC
e1hT7i4iRJX0UcKFseU1ttL1ZJyBr+Zi6g+6Irn+fBorAkB/Xa5baCjd9TWbuBiu5CBYPA/yPBpF
rL2QdfhjqoUu2/kB4hlT0HUtZuW+euS49qmmKTuS8dg3Sv6I8fS5GQEsS81iu2aRYq+dM7szSZbF
4k4uTTb/dKEPvfeAxUQ6vM16+5YclBFZYCO90KyEbH3VmMMqG79bSNysXUoqdFAIKAtPLWsXJGmk
/rvZjp8y/OjWRDwkd1AAFIW7VjeSQ4GpalRJ0p6XIeFbnfjy58kzZsoqfcAk+9uNjmdSglR/NBMM
gUtpE/F8+L1AAn9bZjLy9Pr0BpEooc5mgJAwRkNPPD2+upkXplV9Pl55nBxPwf36LY8yBWwlm9JN
e6+4DLSGIs5LetcnsOKyXpAd1hByCgYDlB4Rk8rb1FiPvGXAtDqGNA+sRAJPPVEs6KfBP9tL0iZ4
6hPKCrHT1b5Rrbk+yh0lMaodYQ0vwS2HPfqVLRrZRyX9Jd5nB1ipiUWsjCjhcoPpcz0NEgx98Bcu
AFfBhjX9Aor/Dnqh1I4TxYKLn9i7vbwq6DeKm9UreS6pc9y+yxIEfdkw98yINAUuIB1aHTACOY5A
Cs5WvToXKfuYNGclKWgQQBVkbGiCp0Igy1y/v/CX1EsbcJpPWqtpBGhxORe0O7QSyVd5clRfT12W
kbiYJ8sCk9+yIbFzkYDrDsW8muggFaOfA0/KQvGCfDYwDSP5w4sgqsm1gfIbh2lSX4mGVScWbDSD
r4vrCLtqt9vY4VVaDrzxwBwkRuh2xhDwML4j2Bk2VX3TXkwSL+VOukyXfWhHY98m7ca2M43I975y
W3FnSm/K5ANPX8iTt/EEyHGERxy+EcfkjAHGzdrACVbxr7m/GUrYQ2TCVAf4XjkE09LZhA8P0hFO
fjmNgbYtaoY2dukxNAaUr2zULmeA9PdPkLAxzQz3H8RVSX35pGe8mPxXws31oCzXxLDfOZXWCwzL
w9wpMb2vapPR7GMd2PUCRj8RvJ6R0InDWTnazAkMYfktU1VT6iS/gRrLe0pFJiVZ2sONw1BhG/Qs
fN0G1d5rq4puSWi+vJrWnFvtyg5IrROsZXckBkHQtfpmx7sO5O/Hb47qHIb/cEAyVhLQGJiuupZ0
PSMevHHL09pgQbs2Sl4UfK/y+WVOXrkcKzVz58ELeoOHZObG/idZFU/wB3nfsPtrwEtMUjdr4Mpo
gKzhdxWWZ3nUaVWirQKbMjMN3bXaBE7qUJLOZygHS77nMBM9BI715QZunujXU/irGKsJ/0QBfprn
15/mRUPGBYJdMjTH+BEQERDKguK8r+s6WpA4rWJNmvW1nHTiwJCYnzjaRljYI+NhL6Z4AHkdpZjQ
YHsjmaxwlOqVb0NArpt6Dd5RyHeIc0XCy5bZe0bcb6izH+XzQT9CIv+CV/nDnSUp2Rgg4BoVaDF5
eB0NQvplfPpsSywWRdpOpkg4Nx0hNNINrT6b3s+F6zSopOSh44BqI0QWmY4y6tGK3MuZs6TsJPh7
LPefznXt+lP2DlG45o0VqKZytgZBitrjq5WvsNnZl9Gll4lhlgJJffT3UfldCCeHZibi1Lb5TWtC
DnFMT+HGJR/y4JcoI/ilhftJ+i1pWyV7qE0PjNbH+td41tGTTIHwm/ja6SXOqDN3lpb9OEf1LovO
xfMOd1Eq6pAZUd+avWFEMj1aCiyNUB6HWA2e5HuXTuO52uOeW2VzdMQEibROMni4g4VW6KSRg+W/
i7EV18y7m7DUXJBMrDWz0OsARe/yWWnDZ5XhAwRP+VCX2EaULKDgR0I3WM2w013wOWhJvBuOljUp
X8JX7adlK4VtNkwuv44Qk+y1x/L+pJwDpySqs/jp5NhJpMlaENTPphzfKDEA3j4sdLXwqPyiNSUG
VL2jMjH/r20QHvBdg7ZUiF8RFO/zBhnW0+o1/vecQE9KMGSbGroKxlYdy+Qabcn1qAe96oYLPyhk
g7t8i/lYaqhhAz9Bh88fd5FMiXD2bXXkZKmorMVBjtFYobFCUIxSzf8jMOi/I528Tffgu5+ldNVe
mnlN4GUbzOu23vTx7SWecHpWYQT/ujxR8FZXrt3EYnwSLBLnYBP9EOLvEDMzqhUrZXnwyQ8RxcsL
yAay3MjtHCHkz3YtRVFTCZPKNY76O5hc4sANASvK3UvsY/Q1EX9uARqyQHDPZX1XhOrSZWzpeu5x
hlbtcUPd5skn/IVFZCh3Oi7EC6VBK9v2oGBKbRimdkqSf1RACfbABOtJ6/X185KHreXwZQaeTot+
RrC3d9jQI+e5NmTS/yUI5AM6sz8P3d7k3LhqcB1fJeLU/E7d5q7dA3LciHbdtyg4EcDXiGZdbYoF
NcAyMxr2eh7+37+1PGWDroM66SocUGKbMkvHE9AorqdxTAhCK2MyTVCWrQX/EhQ+CHaQuzt3+qsi
u+yBO4nLZ1DbFlO5c35QpsHdV6pLXdT2jw8CKvykx8HmK34B7FLN5Fdlj39BbaiRjr+avEYEJEzV
8+syDVEkwGy8BLK6juzzblFGJsmYuS8mEdIZOIKvp5XLatzVW5QVcEcjDNl1WtcpB95966Ckf3er
IGvAzBUCRR5R4Bgs3ewYXqdfnKWUOsJqmNI6L+kE1SoiNPTx3XISLZiFOciXln3+kfElpNQMnd6V
ews9qCTohWmM/U5eYEwRkX9wSLEJ6e+kr42AfZtSFGtYZ9IWzuXADPspiQ45B4sd+MRIG34EenyG
4aCib25LgrMGvSJBVZESa+7d1jDeFEaJfcQVbQsTC8pOnAIwnKZDbQazmhszsNFqciqnA1XjY/bz
iYNaRt+f3jdUR2F3p6r0keOMaXCCQSnp0sQtPGf30+YoBtclBgGsD453bHMUsxXBLGAiIuA44caI
68522e2wblYOASS52XQtFCWlaTp0TzN8esf2xN9K70BinAGvzcpkBgmhw3zWEc+5SRjPV40nh33G
0+BFbJrJF1mfGgho0GJGvgpbnUlfIyMgrdyQfwgxmdDy2FyYTlH5Lh4IXFHP6eaRDb/ItjZovUSU
sYNOZ1XASgPCJpz081ZmCqwVl2fyekhYOSS5SYDRbJzlCN0Vbeatj1tgj14JMYi0tJ0Acc8LqnJu
7BSJjjEq8Dno/px17lvh+qhAq/ELKvMeh9r1PJktc9bLV0Pxyk5m3E11MRTwH5FviSnyD5Pao5uF
tLPcvfN2fP98UNo/55Q1YfowNWIDAHBTcROKUegNLr2YE/IDhaAwTynTWsxCl9WO5ankniHkygVR
xbloevzc7yQ16tR+E7AvYhw13qx4q2hfG1Kzhgc0RL0ikxa/sWju3XEDSdX83pXQVRkjNs+MlViN
SyvneSfNkRpnbDyFneo+ToAksYuenAMqWI0Dc5YNj6LAMGmZjEgm81Rj/M69241s+qwdQySNE5P1
u0gIjFVs6M0U0LWls5DVddDVaSzohL+VlWUhERljQnxCzniUHUSirWYr1tHqFG3LgeN7oHzUWTci
m1Q8u+w/PcuhA7R4uqDK6lhXbbF3oLYlDT/HFISTnR0NK9MRmfPe/vzNNIqygI185faU4mKqPA81
UPkLoApvjXxFgfZrrkKfHipW4gv7ZOHrMwrria3XA4N/CFqX9nTr2ROweW2cRus8Qzr1et8E5Ikb
f4zZWvZ1jbBnhpI3Fwg36us3NHt3hUedpOw8RjDI2DwqpWCzbNOnN6gmyKIv6pkEGWRvmh27EKLq
9T5S4pKfflM5KN6YcONvT/yO7TlPLxNhIVO+ITwxhjALz6xEA/YYrj6iKsDvncP8wFc8ZPQbpeks
/4/Qk38ewGs6wy2irL/osSZA6cwVFouiGJhLRZhIMh3iP07g2ZZDFtVkXeXLizdlT5exYoKYpOmS
4cW7yeowXMS7HhDeyOSxCpjWKPX3LxilRFuCVij8hAj0KFfiNt8tGzRKsVKXgqZCdFPMcvhQrGvB
rD0M+Uc884OMhKthFf1AgvH+ZwM3wXE4R/2zFMu7MElVh+pWZBs49qUUg88Tm42un70JqYZho3pV
MQ2khh33GKZT4ThMjjzbdrEviMk2Km4iq9t1hdvqr+gH66zgT/Vodysb9NoNHr2EiruDDQ94IZ1Z
us7MQ77x3pPyJ3+JAvs010q0P2SqKkiUJOCjh4m7oI17IiYh593sLmspCgXE+6ONOL2sqUhcj7R8
2f7kqhaPtOj5cZqWZDellXG/t5WB9mNqRGzQakXStqDgAN1vQhU87Ct3lLvkVMxTqXCZhTYRyhLZ
Kl7Z/CrbgWNshmGSAqySd/xcLrYiuHPvCb0BpvomF//qcmqQ066u8/8tHBS94xhW1ETgKBI90T5x
zKTVCZdbtSVkQt3E1S+px8M7YwC/5lsxuUAKCZoBVUxAbYN4VU9aMYjD0S4fhZxMfyTIrOhAxTWY
yHYx6CcLFpZT6EdOftlapexBAcav3kQHcCIH/i+xa37z/rkfBV1jrZn69nOQzLOm5V1Ga+xRVFHT
IflA80AtyHJ3nT/zP/GHsMxKMbqztjO8TgR05/jW6al5we1+8ns0ASfHfvMCgrchhmMm6Tr9wy/6
Os5/5y3eJuCwayOXTL/63J5D6bCiLNalOyGpbtmTiX6ja3vlM3hvDpLq2Qrw2Sjwx2Zfmtz4v95G
XmJr2MhLLbGreo70qCs6zV+IjrOXVJ7VvF4dxwZla00F7aQ1WLYn79/4Vk/XNV39iqtR2zrMI/ZT
1URiIYDLcPHQI7j8KqTUkVKQOHVNGwxVp6wgWNZlPI1Vnzv/4lw0TpVKyZ+yTeNhXankP/WnbYkV
1Oj1YoAVDZ13U0K+bQ7fe2s8WTp6NNONgsdHpYs3MmqNsrO0OK4Cf6WrDDjdt1GuIdlTtXUuxjaq
GEHbF3t8rmL5PI7MgC2w3HT/M+A+8TzKXm6sqU4EHOvfvVEgeR74BrkBxzCXmNxIv0UV66uKw+uc
T8tcrvEj+A1axStaNSxNXF44n1txLp1BtQotpEK+MX+eJxR/gezcmOtrnFkIVAnzitRw/3uJGxcP
30H7DlGHZGBT1Eaz9HwPXvfk1OfyPjIH3XH5fQe9uku2KYz6ldWUhGEa+T/ouTilBF9jiJCIm4Ld
ephrR6QcKDSN0QQcfX4Zgz+ZcUfcUI7+3T8gXK7uY89/LbVWGRdiAZOxcNF3j3Cl9C5dkjBSvPjS
6QGR1HFsxPdTkd0UG9vG3fYJxVQ96rUC6k0bcI++MTaTKFNeQlMMAqZBLkqxX19LlVt/dVB5QBLh
ie/LhcbhBdVdrv2rwevSOIlsu5bj+J+prpteutn0jfjVXbvRWS09lKfAt63aCUCd9CsWVpNGe1Fr
T2Ajh8l0AT91gAQfSjKJjibQuup8lum+VCb6cKMwFiVVi4J/N7Mk7sFgBoHpvM0NMKrpZh0SBQ4s
ag9VjxYRqa0gB0vjfgoAW/kKdB7aH4kbxQefVEseddLvh5eWT1mPhQioqpW1WXeCSi4Q+9jQ7mZg
nfUA9VbrND3KD230mfhsZV3ztqvpin/ytJxwsjoPsX2IrjFjTi2zQaTj932P6saBeZktNVQ/hT5v
N/czspyqKWb73XgJZJmQpmkOt2j1qHpve6L12W+WIk+tF3F4OUaCUIDtbIGZaLx0mIetiiY7wiEY
eFDrH0CDDLrTKmFSYy1m8cUoFrON240GuPqdoDYqYrfpIG570I+i2InWFl9+4hA0hCsXECgC7WLn
O0lX3b2eVsa9hSMNn2VPJfz/UKRHG8KTUT9AeSHfwYqc1GwCM4N36cFwYToB4mo7QFCrkWgslo3U
UM6+8JY4oOsfgBTUbsVm2msJCALcr36fechFLh4PMgzSQD9HwFQdvgH3z+zhoRbrBCIeT9CWxEzt
gDFQlKlHfpbHhEn4CGXOvz/HORxdPo+9QMQdC23Qp1/qrkh2K3ZrXdgjh+8Jy6U5BhL8cZuaC08U
jbfKA7AfkNTk2LxJTfw1FotCumhTsr4wjODWrFpE+5VZ5NFF1NXZoAtXgdwhwxmNYFz9Vmqe1Jk5
xFJOrE5LeUg55ksgNHsAm2XRLJF9VPWrlR0jb1bqzjQ0jpb7BoC3ioc06KjyWS0bR2P4rktf0J4Y
YXo9qCW97LbkIvsX5ABjWR5cvxrOGlsciA4SID0O8HbeehXlXP0teDi2dzCgZlotxVNPMCljoP06
hX1SxKW/gNElCm8c9eizaI84cV2Y49BwLYdNz28bl4snRHZeuSzf79g1T6c3mmDPt8TCwNFtlNFY
IARigaVbAHqkvAWechrEkqxsKQEqmX2IpjVkAwchxUWufna3gtwvk/bHVPLpu6ReJKb6mGwURPwg
orYIqntRG1FDLSJbR388mEuo2myP8bgv3lx0YsDhV6mTdxdONZYTjj3+hNNdP92vDxtD3PfeHZ7O
bBlh/YEg0YgZWO+qXchXurnjspD2nzaHMzQbDMkAc1E3sK3rou5NbQzViwbHQ7KXd1JkArBVPv+c
+zA0jFQUvaZbGthb/4cbQHZV9+suVys6mVMFVbbv/eEyCBmsozxqwpSwV/iktHp9GKuN9QWH5l8n
8OptQQ3BQV58k/E5g/WqzhJPKu/CUTZ/F6KJn5MAp1+dkC5TLC+LOvyF5A3l5f+0EMaHXrV+Xlpz
ujEylZWia67KwChY0dzyepFuXHn9vBplep1DyvSlwWVR+gUnEOe3sVPeSnji97uFoXEisS1IKJbK
M6LMq1b4n/mJyxzsvf3De2R7ouQWcrCqnyTrc9GIens6SzZsViG3l321KylCYg7DayQPNXeznTi5
kEtAoTU35ABdM0rm62/KSlI5Htorxp7ikIWHlYawkdvz2s7BvQL0tR62r1wrmSURnbv/IfUx0PJx
2Xbz/rshpd4nVZrShZtUYu18Ti0Z3ombaThgwZO0EkJqXa5joBo8ABVohAOtUwfpDdpmVnBFBltq
lInLkrqFbqspzlGuE/0iYNWac+XjCDnfVhUnPE/F75iKF80Wt+d5tyqHqd252d2SgqSuujP1DDUi
vEjFkPma+8nAHLvKL938P9836G6NsSTxs9e2+I5tGNIVBLu6V6LflAS5Rs/jrsIcdWQJ5H6R2H2o
N+WdePSnEWUQcGne8VtbqNNU0XtLafvUy91ZyQtTdX7Su0eYdPyx73NUO8VjBHvogDvrZ/JhssMW
2LjAfFMCoMOyj9terGSLLaFrxi1Bd0NiLZrOu9fw2DW+Tz6rzDagfks8exr9t7qr52vPXbQfkUsy
e7Jl4b5gF1fldeFhln46QTSFDRAFNfCF7AGgM4ddpOmwnLMSLNb2k6CkQFS/h2lhdeeKnfOqA6KU
tzgQgz5XwFuu51DnZVeYqrZnj24TCm/W36GAb3qwH8wxL595ArmuFgaWLN0ew8DvgzPVZH62OeD3
USE4IoBIthdWah3MsrNr8h7eKnz0bHBjqQJgw/ZdJB3LxRrbjG5OcA0KAnP6MuboODRM/DPM8yG+
SSWyc10y/hOBPSvWz/Mh/BxGPzQY+4GZiGVT7sYB1LpXQB7HItpRlH6W8OMlE5/KaEoF+IeLKUKu
lSo+sGxvOTLzC/URFRYdeRJmCC67JlPeTbx0/5ol592hA1RY5TsYnFiHGucwhc8Xxtnotd5ACp5W
6OvXcLaQFEqSRJiMfnhozJbfyS/s8CaqVZZ+cY5vALFudOacZ9bIrkfHZKWH8AswmghawnFMqFCE
6qwZgwoQQevWCijgBo8E1nk6ZlTJKZTcdyDCOucg/RiC6biue7iO6eOoccja0pE5ttmCxArmsgB1
Q8VKeeRchyFEL7GEgwFe6T7LHNQiVwcyvqw7bmSfI5OD5u9mXOALmPOPueZm8hZKwuhWsJwkQEqn
bxkbRIpIaEVg/KK1HSbT3VEv/FP5tzzCwlnBnB2Bs/50O21xlS9aDbWl4dSJBpb+GZdPO9TQ4weZ
oQddl2X8U3Bum25WIbx1uActRADsRr405GoNlW5YnH5jdQTkXtn7o2CaNFMgtYKOXb5A0Rr3HE6A
4OKA9lKOM8NMiF57QAVNSyMKasrbCE9rQRTf2RIz+ZBMpSwRTjbvs8GiYoDU+sZpmvPjpmVF8h+x
opp9j9sE8Eu5q+KYbn455zx6B4NqGGzfksQSGb2rjWnNiG7BuQN9eT6oBGQkMcyu6Fo1fWJLUYlI
VEZDn0MT3WTXFcJKccyaDyeceiRQb9uT3/CRB/zvdjdTkH0ZuYs++WF+ok5jvgcOs2QK+KT5qdQE
17akHTgP+ATj9UnmVg8r4DR9tEEqwNZds+liFo9i4a3I+jFYFUIs3OWifwOXX4Xtsnpu2lXPSjij
wa00/qrfI7V63UQZIvvJ3I1EN7G+kwA3Xw1xN3/CLFKCeVAL4Y3LX0Uy2aiRret6OwhGxHCvBWL6
8vd5Qds7KgPaYnbVS2rQ7RRarm0rN74sRJt+hEiYqdefFDZW+Ayy4Aou0KYQB52Nyr56z3ZJ5wEJ
k2NWS6Ir1LqnRfX+SDEtRcOrUttP+RCIVp9/DDe68qPwFuVmkxIgvNShsK2CKPIapgbKLSGOyvs6
8peZCd9qHXo7x/8MuQ0nDmNTlX4HRuazNnVYo2igt2k9rviqLI39EPzRV14hYxWsUm1ueUN8rIqU
qlTBQmndzu7OWZX/Qp5TlZowRtWi9N/oQme0WB0FbuxLgJ5/Q/LknU7viR4q3x52H2mnk8vVcipR
ZZ9HmF8GVM0DodyjvpWxQ7zJlZ9C7jtVUuoX/n70OISHePRq4n/uT2203o0I7gM5gosj2g+P4X5p
LdGl8EVQULxam5KEp0SQmCRGrM4Upn4tE/I9Fdal5iN/d7x+3HWtXBsnljHwHAAswsCb5eAmMc1k
CFxAON+I7BODmG1f9HSRp/SsjeqY2rSS5msai2W496QieQmZJrAdxX/aqqEeWVeTjOvjXf9LxhQr
Bt+i3fWZ4+bxLsQ1NwALuSFHHEAIOdK/Na8T09XiLKH6b7JdA0gJLXOwKZ/jnNePdkgTKa1j6tZH
0AL+31g4DgO2glA6UPb8ad5iRJ64wRZONP6AZMZX58/ZX67oRgLcW2YQH3pnfuPk4pqMObrQibVk
R7gwR7A4Z1rAOO+LPsJODA0OoaBRqEQM20y1jwEIObz8SmYf6nfphwAgpwFba3bwBU1PHFCmP77F
3WFlfSMXM0dJpOrIWE9Yem0rR72ic5p5q4yxOCRvW1+O5V3TZ4z1gjHAMSZxcd3fF48ilUcIZGFX
Jz2/yM5OQj/+oYWaYiJDhzwhzisUZByDbq2Ibs5m4r0DC2L4zHytS4TmO8Ifz8ZKcsu7SZ9vnaDK
XN5I1iK6QETVwxwwNLcOaQQVsCA1JASJwAe7uHCRb1ZgB19yO6AUEPqsiwYFklmFeWsUDyz+6LpG
pXaepz2D8EgZd34gL489eUXJsvlS+bRzVGHLPX4kId04lcEsHO4s+VGuQapDsdMAfEQ2Rr+iQju0
Z4lkcGXUEL4do0wlIjnt2H9Un+k92jXy/+fHpAxy7uLILStjC9VqinKLwBDSrD9eEaGHss5jfOCo
O4qdS6I66aviICfAegNzSYHiOumX2bjXiUM8RCAJmEJt+EolFuIO6YB8RElxJLALrboFVF0wOvUh
9tV7MXKgv+h7K+mAzx6tD5b92iUu9VZuY+oPs6uHLJFJ1wicg3sCTGhyqViHJNHw6sGiGdWSAsTr
3OTMXvv5xMLQvnZvZQX0Gh3v5eu0sg8NV8coVdlJBY9UwVjm7d/1IlzvNxZElYA/Yc3gGZB48Kgf
icW35LR074J4VRyrZCoP+6Fj2jmdYret7ownxyWygtNPBdXvzuJve6GuCYGjvfhrKmwxfPkEQbLw
MJ70ulBChmfsX7hJR6xQTgwdI23I16eFFaLwaAt+KZ4w6+DUYk7Vwyj58CxOWEwhIm5Eilz8mpQ5
0o1cfmRypoibBqViAqLWRU1PcMC5Vo0UPer7l+RlLcUJEmxQWX2FgxrloVfY3gJy4FVn61OM4LfB
TqBLTCIv1EfXE1+YM+Si0eqmPBX2Pip98KNxY0ejN5QZfY3utifBNySmbtJ4lWYbWtbtNs46JZvb
G4ybq+N3uOS4nkTbGkOBgg3JxUdJcRrT2fqlQVSeYnV9hhSyLuLzSB2LYucFS+4Nnr4WGKLN7rrg
yCQsF9+HSKpbx+81VSxlDNJAcycizKFv7zXSybtwZ6vjgQw9DyZKNIOYGOgYLbnfcZh7wUjsnlBC
NTfGBlDI9LYsgci94buPlWWb/wi2kwxGyTXXTTvkEJPHxH/5chzCB1TJr/dYWMh2JU48p8xp3xan
vaRi28nxVc7nStEoow9cua8EFlUi+uGT7wvb4/H9aQnhCT05+56VuoKYpgCiCT6EhBm4OfUuxZrp
WFNQoIo17oQg48mlhDi/lww+2tvEBl3jTvevw1tP6Yk30AnRNV64ptoTA5VpC0oRQJOk8HYT+ofP
vWVvoHT+EdxYvqmBZHiuGvBurQm0UhsvvkSJr5MjgBeymOprsd/JoxK/ra7ve8Sh85GwjAt18wq1
ckA83ySuIv+kPWz5BcFFWNSZQvmINak4WMwcfmlipSOJrJrhO1UHVaozTyN0Gn71gPVs6knnnpbF
HRCHbJXMTibh99FUVuIPxIzYOD5B5j3YVRgFwBRPFT+LTIPc+tAe1Z/oPHolyw+dkMuXOY5QTX2T
+u+DmZxLFMZiV3hTdJlgoB0eEJQOCEDv231maxqGQn0G0BL1Ycl7DV4g74Q2lUKS4E/I78lqRpwe
DgWOzybWfrqb9iiyX3fgCp8d8VAv302UuRBuGnLTEe8kl2rLcE2rBw/uOF32ZQuM2+6isqUQaSgZ
itPHHcYovYfehHdb8eUwK0IY4xSy5BTHzbTbtO+YXxfnYa2WDc7nft8Fy3brxQK20FgeBAKKlRCt
1bQY/yDGjYmuvN4B/UhkTNPRE2KHLKzzhK2C7lg0511GjS1a6TnC9fLzwFN9uqicVckBrFV0OmkJ
YJLC47iS28juxJBeSbhA/qIcmt/ZGDgOeEvY5nAvAuKLDfmin4I26ed+CNMT25UeTXoXFplr/vCd
tXquSX/xngmXE2Jci4Ee21SL5Zf4mPu6XmaJL3ThMM4uW/umMiAN9djVZa3EzenPeR43BuDweLB5
vaKPQAiepytvsekbrtp2JTkEzp8QYD0+srEa3rn2xyfvkWPHX0mWwFKDIujFgaTrORku74gWp5MJ
iVsBg+7JqFj05eGqwEBAESZgQJ4UM61kz0XPqMFhhvcsf0GnIopxQcUvyYNK8T7/2imtS6ar/OMW
44QTNIURgQwpBOXU9o0FPFePsbdeTGQGZWuLsfqVNwhbBq+JoHB4awSFk9ObTXGrgiRDKY2PGj1H
ybh271eyA2Tex42h//bPG8Pxd3uBkwBWJ2qFG0rNc7mn39ZDCKjKVD75m+lxTCHH6o/8k+ANzH4v
sQwi29K5dytHmHAts3LMjBbHZAqSwZ6VHpY6cKYL7wxhlblgES9aG5KX56/Yn1jnojNe4u8Niux6
ig6ekcsP7lzt/tuI7We2kxcqDtLE2C4xqt2AyjEVBUF3ib+FNamuiSH800RJiMEmFkBmHY1jsS2+
4T5TbnNP70jHsZOyWFgcf1Ptl8mz9QaG/eMuSUDWBh+9GZQYCz1VzvDhAIIGjBe588su6FBY4tox
/NiLbEtBX4wKL5mbuBSNqjKlAkVGcFfqTXBrL9HgQC26jhhWSQbQYltY5i8Hzwy1gX2zYLxo0gMF
1QgPmu6nOjvC+oDxjtvV+45jBvn2fIDPrQi+3oq8LYytqOkICaNxpmNRkfQHHvFDD5uuGB4ffur2
TbMazGJJgprW3IpH3un/iieJjwNhuQenI8XySwsQ6o1w/BhFXpYlOjJsn2l/4D9NzuOPDFY6ikEf
fJqnSYH7IUq1dC4XwRtoQx3QNsVjownBabYxWmcD78zfTJqAxkkZL31H4YPmb3aLtnJ1PaMlvaGv
Vlw1nZYmZokywla3udVhGZBVK0Tr56vMzjxYESFUKJHCmvC3R1Hx1GZGc1iBg6W5IOcg3O3e6t/A
hi7rzpWeqaaWFQa9Hhy/1OnHtt123MWkgHPBJhtcdGSRorMGey9FYAjn2UnbllZGd9/gK0lIGsO4
WsQYU1X167B74Sz3cbIVHMJVucm+segKdSwmV61gPID9awj+XxHsEdk+fvk4VScn5BXZDZbL4AVb
5dRt5qfYhpHa64xOGEOwMPp++ijMqRPl9483gzfkYtGsZgBUOuGHrBPDTErm2HQziujpacCJKcpi
pOVtiYaV6eMrfX2Em0Ii5ihyyeLyWUTin+LeuYTcbu1iI8/I8kFqB4McAVgMV9jV9UtxFc53ZFi6
GX7bguXyg7vNAW6huYRAeHOQDSS524Kqa+ZR9xx2hogiRbDe8aRlX3uLJwOJ5wqVGFzJdesDoGJh
+F+5j7it7XetHD+/XsZJKeQhpK70XqCeniU0/WEAV0SSF1vyrmyqqyNBC59TskHygDBpxgj6SRJ8
dwtAZKxryPz72Qfewl+gc0NlsPigvWfT03P4p5OQr09xZohXixKJIieCK7B6n1On9iDB67opO/uM
uLWeW0dIMswEPamyJnkJ6+9bX2F1o7dg9meJn1hY78w6tiHXm9Y/VG3sfy5Eqx3uCxWEOe87+eqK
9pwKpDOW+stGzZxc2wUgSUwFEkqFPkvr5a2bz8/OYdExOZecRekr5M9d1qMSRZSLAFBWSgc/kPjL
uKvgg5ni/aILn9GRrvCkeQQjYCDyQWmn3f+bcJf0SkpUFUnLz5+upfeTbWv35RutvajWJyf9Kcvu
/3h8wxanksyVq3EIDJ8yxgPXc851tw7a88hYUvVz04O+Sdp8FXfCnPvRwP1hVbArxW69/NaVwxuB
UGpAGdOdlmu4rv5/WZplAhJLg1q3eRUCYX0AwG5sjw/LvQwy4e8GjW8zZW7hP58LDn/+hEuq1io3
5Ws7FGcG9k7/6xwjvxTvpCvktziftzYumLQKbtfb4R657kMkoCb1LKYNkQoqrnLv9g9tpmXykKbW
LHQ/EI2Q0KkeNzcjP/mDQQI9+YNkca+Q/T/Gf3y3iB1G/mekoMekHFFuiy/uXvWnUCS2rSRVAlhS
N7XcvblkoatNfkAYnkhPYBM4b0krlTF7Qr7zZFIu+xbonV9TQFo/i216zb82qX4U7/OlrHGCDg1Y
/0IqsS9u78eKm5Up/DQ1CvlQtO43BDeBcj4tw+5iMY7Rlsyvfat4zdKlAXyHpRUsRSqmY0n4uwQS
/1B+eI/Sf3Aq1IynIFvyezTnCSbBoJlRochAejx57ataaw3ZiqfSgYROVhFzIOg/VC8y1hPAxm8g
fNTsMxEqCyhgoRFd6Spg1rEYqbMj7guFnCOPE2Jm+2i4ZARjQOOmgJskUm/typ04FndgkBhES0R3
zf26my+NWVmQ6M4crMqyKe6hq3RgAFHvf6uqx8ih3V7NpTlbeeXtKmo2+qKLhwvMr0e7VbOsm1zy
lgZsofTvrQwK2BQmwrZDpOYNWxqccl9yNWX5fH9khptllZMb4v3YEPtYJ2f5vzY8b4HlwFgCNHGE
83Sml7PHMYfCOMk8uykswNd/K6F6SDESPjf9yXb+lHDBuX+2a6HDhpDaVytiY3k1w3wljX181aC3
Wa1xzZzbm9ySdPANJGEsqcJbfNBKMJoKHdNJIKNt/bs6Glen2+R4ONMiHG5DGnktyUucf9XnZfpV
b7Xaay3nNANTGfkik5BseUOz26RnIdEbwO5i4ocy7rJy9lnqPNN7IR9qzeLxsC4KuaGVWXI2fykP
2faKKnjNN7/0R3e/1ZBgCGqVQOkVdZsi1+F63wWak0LzqKlf9XbIosVO+YFVWm/d8LoOdYc9GjyR
ldvheyWSfHb8SoGQ8rtXEJU7GVWurpJGBLBIFmAbMVlnB5fwC8Z4ZDCirZ45H+gtH0Ujmy8uggyi
QSZYthmypCr3MX7wz9mJ6fnKkyVJreW8pP16+ISfty29ygZ3jlgJ1oCGEmrWA/gctCQCK48FbTZx
JkNk0GxKissjejB+XdHG4W73YLmuEFHa5zobu5CRFYNDeXXHQ3OhO8TS58SF19Y6YpWHjn2mFc+k
SvYBgNWa+KIyEjqyrAAraxsX2glqC6VcY77XTRUlX6WYeNP/FAwaaS1A9voHfZ+yd7YzR7ZyKBK9
zVYVqAhoNd2RmOe2MYTmOOksTSsF+VjyGvvO5tCzai5ZouNKlxSDcWJurHTl3RHVCK2kKhCYAy8g
wn1s8W3bpo5bopbBMwlPov7RpB/uz7l2bWN1EiNy1m14RmhxL2z4/SHhb6hRhgeqenyN0V55Yyj0
GDotB1ZsGuqQaPhbs6ujc3yVTNmyibVQF2avURpCI/EJaJRyiOd+iPRjCERb/2SDet8Iu0Ix6Bev
RKckI1yJ7mVAmpY4vcPpZxqSebBSS4/1uQeT5BYzFzWCrzp1wJvcnDoYV0IDb8QtiCzYinBWDsbW
BXkuSMLfTyVh4B0iYVqDug/C9x1cwnVEU6teeK6jYHxhY9SdU0kYwSZG0yASSuzOZbWA3I9RXmJ/
wn/q5ebZ3gMdocG9WYNRwwQ8JhNzgm1UCFDx0K8jCUoMZSzytwmY/3a+BxA62Fc1CuCSoeFidRzC
e9kIkx6m6HOpCZQAe7mODS42mtG/ByxLjz2t2N8xdt1ae27H5I15tGibBoN3OsESb1NrIuLa0E4D
1Y6Vad/1PSmV1qhu9dRt4pLJ6DE0LvV12is2PxDL1kI92CnYhZKO3pwr2FM2VZ6vb14ckYzk/TrG
T6svHMmxf2u9R2sIwv0/DQUhuFqDFVv+gO/AXRQ8lYvS0JN/Naj7tOF8B5ebsds91GniOoVWMAs9
ImayGSw1zMj+kqx87EWOpH5R8WaNCLMQ4MVyOvUySBiyAynDdJ4OyhnrewPhZXE0whgF/dWlFnN9
CewmCFNl8cz4oLLxPnMzYWhUhTYfdWkase7u1wjTib13bMMMgecKS+Nanc62LUe2HELCrFdFZF23
7PrhlhvajnBIv2+raM7neaE6hLYHpOJnp8OMknIUEoPPB4O5AU1incfSeonvrrUAcIjmzmu0U1WK
jAe+jjagHIrpJRl/sNNSOGSC8E7Ypf3Oiigqp5d/P6rB4y1v+DXDms0t02Q1rQw730n+vpWs299A
uaS8OWBlFZwVbqPTI8OktVbJVmc5kVFe5nCr7apdO6LhhsfIjL1ssNddLNKJSsLRYvpcVIxgX0oq
S9orqEmdhiN7FCGxWUgsGGPxyTot/EmN420SJKZ3uFfAxPkr+7njNt/S6K9ONLEikzoMprWFg1iG
L08Bz4MuXX1njOzPKdyEN18SZXzVEVft85UjWLzlgvKy804zaSVBEg+ExmC5lZd83FQckIktvW32
9aYoXCfbhdR60QXNJ258LP6GRhpX04MAnndFh2J27fJTUbxn9q4C17gIhjWAIXs5u1bvWWY6hNoD
HKR31QduB4yyVRCmOkOPBNALNtfcxMcXXXWfPcMXg7IlV3xndd6HD/RjcVIyQzOmdlrSyENbgdzf
ywrGVMbsqyYL8eIxHxFhWs51UY2cZST3mSXfPAdl7nkGjIAqn/Aq9kSFvcLLAlW3JRQM/PsXu8Dq
cgYZPYBjoI6ogPaaSHZtoM8Slz9qSrUf8admguXCly7mWL1zxUTimR/X8gpks6ivnkoua1Bm5uC/
ASw1nv6iY0IxtfAhh6N8fVXOUr3wGtIFRdk01IX2yM9NdjRb4yaCL2T8KGQedJdKaYQCKhmxBJSv
Y+25UJx5mzlBa9vh0F3l+pvk2CCdWExKZtgDnZbzIL5Rdb7DEFEA2/VZyKo4ED0kMjE0jCyW5rTJ
zs7C0c7eekQLDvuStvuYlNdPTPvwwchevKDrfOoFCnmF0Ev/lUJVUgXmkwHIAs57F/X9ffqi5zxb
I9/KTkjZnztj6V59eLNRBgKqo/jluw3/72DqpIpeNQvLe7plkXj52TPxaU7Cm2K/YNXO/T42qiBq
YiWW0V2rfyxhqobZfjmk+8japzQA5/zYpWCFuUM42f3djUn5JlbdcAxyLtZvFpMkBkx3QPdFf31L
pqvPThisAQERWlXfp6jDdhwwfbovJQSX5Hec7G3ZO1FFZA3Ye98Fu89y1BfexF8x2T8dRuOCGrkT
w+AsJBsJ3fHYiZ1U/h+sevOehZUeK3xTAnhBVj4VcTv/U44F7hVlDU8AxCDHveahZR6qTVcTlWjO
E4pTC4Z/MXLaCDt8V3YmxPJIvQB2IUoEF/rNdJYpO7LywV9jJ6OhcsHqlFRkhgjpcMoTZ7KvCARB
IABE+6Oxu3ikeQF5y7YtzR7Is0+2Wh3l41n1VIFtLIZ4OFih/Z2Ag3z4wrcbtpOu33rdk3o4Eemn
mYiBXLEuLB6pgssXhJZP2QBKerEwxaCw0ICnm4P7mwHIz0HI8H1CwdkQAMn0xxdIg5lvobGW7ZMS
AJEMkxZlVQ1UxO4uVVSgya3S+UsLJ0Vm8bigQ7sbG9lhZyPL0uvqbCb6Mm0qcD28jgloVovfbH0f
gPcXxv2QQDxKEKGq9b77nc2wRdoqA+5KjyV2am2TEcWpdxhEY79dBi29L3Os5XSON78678lA9yKP
IO0V5Rx+nYAk7tOp+/9DR0JnRGFWiR3CUdubyCJok/QwTKcyER4CyY30Wtt+fYrwebKrpQbXqeni
n7VyiN0IeKg8XZswRqj0mSmxjmw/A77UFHXPSc3z4aHq+MfMjgGiHVkUpjSSU67yPqJiDG/GFlXj
BJ3Rx0g3+HmKP8q6QsrTRyL7KNBB6bWiLb+AE15Pm1tvkA6EbV1N2OMhroJryt915h8gnHsO6Wm9
LK/BtCGtcIqVG5QVTgdEIWMfcMe/Kl53sAJUsCawvskd5B1ZXlT09oGs7sJQnCVt7sZzF/Fe5TDD
bYtFWevNhXEBIR/UvKNIMGMfacIxr9ZrT4gTA2duNc4On3MgB796nMFGodJOB0a7NI97Gzg5uVqY
cXzRy1J8TwEx76P+ZdWKrSP4gWdFD6bZvYuFtc/TkR0zWYzeHeUqrghFvVfI+E3m8YrvMX4Rni8C
m+zMTLBXJ5UoVvXfYgrLSpd81z1MBdwgQbeNqU61TE4tnxpTn92pBfFySuIgr8M1FZtM75f4N8Qb
rcz4+IqMACESkPCoeN+BAbNrIlXIlvs3RWIGC9bMwOtJ3K9sJDkGr5xjJrQ/cmwOFCTmIpxOtg7V
HE36Y3GDfvXPbmtPN02MvUEA/SzOJXwtfQnIPfyg3eL+X62HdYTFFarPj9qEe0aRDNO5x3nJIdKg
XpWfOWeep1p+0IMrcGEWGgXnNAi3nU2QabTePsi95sp5doIt4kaZIHIzOiawA0rrl7it4ZuwAyNo
pOKL/J8BkZv15fRGcITNZZ9K9E2sUQNps2lWlY660gpZvddRt4L1OhRe0tTsz26gps9/Ia7aSVi7
SOVlsbnUOefa2Hide7QmtUH13VEZ0KFFjnZ4nZ6qqB5jKprm2zBcrzuy7ARXOaFXrID5GhdDhvzG
K1hxeMl7jVk2x/980CuZi2OwVtNegq0ziA7Y8VFnXKDhmFDtphPsIF3eYywRjEUFO0fXNjCASJ5W
cveLuIZcAGc5zJ9Dv6VCyiM3coKUAoJ/2D4cwU0OqEFIZExV9V8QlRcS3v/2BJAxTP2ePowF7mn+
5XYrCCc0lyotbQm8sfgEQAMJTibhLVttBWPdC0vPvYvw1d5sFhzv0F8H7FwI/RWbCigfjGQP4W1S
Q+CY4w+D2KG6fM7SSyAaCsQJnlCpwHW3JI0SebCbr/gi8s4SQACMuEgOeBE70yZyNknretQvFLYr
5XHd99SrL4O6yeXikjBqyXdiiW4weTCv1LUV66eijDIfXp8CY9S3tXrOy5iAf1SDPPUkHGNje17z
RwYLQcxcUOBfZwXVzkNf33H2g2Iurqaz3dvogSK8eojvNz/ywW8Ou144BuvXbjHWK+Dd+Fv/7Gvm
BhNc5Z4oPhCsf9JRBWbeMS0kZv04YIwGMj+QJGdg5dYiOOw1H1BqkObs6WK47HOnZ+HvbR1c182M
yNFKxoOpsKYpCvIHaDXahjBe7r9gQcvuJ0pcnGiYQwx0vVBdND1YsslwG14a0RjWpS2LoJac3Vdv
TXX0e/dMHEyMcHnM0R3e/ABgOzSOxRcvs4jWROj/H/6uWleU7/IjvPe0ZHuPhFkJPLXFt9gIfJLN
3uCzsYK+VnIShb2IvSaV9X55TeqszuI8E/QVKc9IgRTomvJMKHNjvc3/Z3rpsAuqjWGbiG+DIjzz
CYbWlLNharaGlugmv/IFi7hKtMS+khCIz70CERTCy4Q/BeT81aVR+raqV5klX2rZ6ePW5Ch9t16r
/393rCMFf3OBJLl/ty6dcQBz/ymKi0kzPTUs8Sm7Jc+5VlcowLviaDjtOMXsqsvk3DEHTPETIhUT
RanMahEGhQTAEU5/OXorCKbpHokTzTgG61ozlfRrSwhJ/aPJ9jRSba1+IAEQITjr7K6Ej0HURQmt
A4lGVE6JSszSf4Uqn1d/HGFAWkvDyuPkR23+YzX5RK1y5nM2USzqefXd2Blf9VUuAdg40CE3HQlb
FNO1r/QgPK3aUbxOv0tv/VotDLXZGjpuDzEPlW6CWWVFbS2c1uuGEq4aeusjNpsS7BTtoqwKPBTC
g8svmQHMxFLotIqYf2O9ECSL/tY0d3qoFJS6zrXw/dtJ6+M9LK9BFRDXMUIgyhj1dhYIXjKxC7cx
OVCfrkZgL2ZHnv9BL2c4AgJ/vEy257wkodOsBy8Tt6ldsZDBIZbiHravUvWws2F0Iwi6qRtMCJJz
PEsqMNhvjIGi+U3ROcDhSTRsuwTkN4mxb/Rk5W4slmQKzujSqTX0cxMSaEvRfnCPROKkFCk2khTa
vo6y3ztMCQSg5LD+v6JHl2MY2ZpfNR+avJKTIa+BNik5C/l7rZ/dq5SKqxCyxpUcbG0a9pAqfl26
xv5IdlBV6UYKerrs05r7UOkiH6USgVez2kdg56ul/KTMjKYqUOiKPiKDFXoqO18ap1JfjgWPStgw
rZ3IqQVi6pqm2FbzADz5MI162CgnHtT93dGwvIHec20g1YyqOdQwkw7FYXfIdXk8P7D92SmDAOeg
XQaN8dC/etnB/WFsC3/mvhCE1YalkQCnbzb88OH2iuomPx10FHYe2w87e+EmnPQ9vqjngjQqZJsC
1RbHQ2+C3dTLc0umoyskJNG4ufmFqzTwobIPaAebvFKdHqNhVVGYAbY904CBf/YLHOlyRANMy4fK
Nvo09pfv8XlwQWUenAkQUG0Q6SufgtNBC5NvnECXyqca0Ir93TUICK9dxqoRcR3UrYfMM/0S3gpO
lPjj8Cd5+zAjKm81x5r6dUsPvEdBj1ILj80wZvlI0vzgcehC0PL4pamW0rDhyBuSszfzpmAJRHDA
e+PN+whdsPdz9ESHrJjDAuXqZ7yGJencA0jQJu4gLUTmQ0sDu6zoW5wfBgn/3DNUcnKEijsgb1EZ
rpUnxIodkgqY0N5oUbUoipHhU6qVD+Cq4jCNEqLnHcQ6MwQ5oWSsO0hb91vL83Cqm8wAstfCkJ7c
lsKZ7DsGMOKTpzt26ie5xrCNCo6Vb2dEuGiNpPHJvAU8uNic9shE1HWt28Y4tpkEek1h+lKagTux
fTgJQ0s1D+y85nrEuRpLNhrzJN1bOGW/IHOd+KrCO/fH4q5NLhg5Jzkbgzq2KJAA2hRskWX6OSge
/yeOrwVAHTLcHnUkSlogc/PZljW7ftg08fO65eQ9gBq8gdbJbmfvfqxw4e2s+6pM9hOgHpFm5yqD
/uol/IWRwslTZ1laLSo6Je5ElVhdEXAmQn67WgsODBV17X/gzSOFHIuDBHOFTQI/H6kdT+x0p42e
qIsY53zoKfzXKAP9Bv+37nYC5wnu3NyVwfmxlPzTBCpe707SFwYnpUjJUb4AICidmMGTzenD2vw2
pYE8eoiu1Ksrojl8N8M5HJdrad0i4MayAE2O61nhZ20QECKSQVMZyOYcral6jDnmqnrJnBCbDAvz
F4qpuem44ZmdlI6WGWsFJp3dZxwO23EaCuSao0eBEgX498tIz0wNLzSLhQMjXh4vDBVLVg2i1pl+
4ifFXVTLuoB1SF5A4krRSpm3H/cSqE4eJ1sbhPaF/Naln8KqZ4rwXP37DBxRsSDsYvvOMxhEcVrR
x29HwWbF4iLGxVu1/KUmv+yoTwrY9zkOgD7aLSyXlzziWO3/EiHr+S6/lLet63YGtET9PHGsVLnc
ZJ32genYh7qQd8Qfcklk29dGebhEkgFkMrwvoxhKTcygU+X3m1MVNGjg6fwvGiUSSCp/8vhoMo2N
d0qIXgXNRg5oBXZO+MfEBbNaibnICfdzR+S3y2brdWVB/QJzk+xp1KSXF1g7ZiEoz4RDgBdblUsr
HoGm3ii+bPEPZR27kK8qe9BnkbRsZcdnh+hrbNxvdRkdKLEmQ6byjgVouNX9PV6ArIJIYSrzcJSH
7xDA+cjDlhkc4xjiW5+6bNkUCD+gyHTZDy0u5dZgB+Ypnar7VQh+gVPArx4YeJhoRPex6RqfSGHQ
pAj6/R0OSJftwZsj998sq/tXJudazHzOl3iSUiuHaeUPiv2BZf5Ggdn9P3+NHOUY23aZkHscfVrW
LjiFaWBbWKO5lgPmH9Up9vbtRkBw29HKYBfh6n9riNSM1747voJm3SSUvO+Z13y8AoCd5Fmp35zZ
ch+AgmUvhEODbpRmokkp70vKZlNCfhpVosQLGqBx0suGlheezOdxk5YM1hcavYyvUOOfzpXE4bgs
DjheYI1Sboj/EEvn/UwNjHGWAzfCpNUH/5r/WojP6KB9GedzvDlqnSrTqvU6BMykQgtdteO6FjLF
0eMplWK3WicQ9jS72V8nFxCn6P60x3YL+81+W9OUPlfU1uoZ9PeTsEqV3hiS5CoUHYHBeAO9eUUH
WT4H123nJC2humz6bwxcqwSQIAvNooZdYjSXfCAcU1PhXUITkgD/UNJzYhBM+1xIce1Fct9Tb3x4
OCbLoB/RViGAiQgE3ZGHKfq6yvdo0fV4pfmuYuYJZ210w6ztC7HxOEThaqSWKByYoovHOJbYsxES
OXTf4cHh3tINy1WOLFCCCuVn1S9J0urcZZmrh88eAkOfuM2fc/Dwx/dHbZz3TODMcFQzb3R7DV3r
HqP9hD4IQVjLANgQT8vJ+dm7KB/7tSHo4mAZoo41WYmBCCEwiS9piW76qGN1VC3EOvNw0RJ/bKN9
6/S58i2J4kMPOn+430nFaVmwQOXPTCuyJTaTySbuRpwsrnvte3L38q2TItuWzD1kXH3ePwylslpZ
a4Xkk2AGqfX57homGj0RTBI5RMxcjgWT05zXVNIt1tEEqUUJPKh1wwuqVidcghi4dski3I8ZDM1t
Wg2CbOEgvFreUGr4M/xdZyMmQsnPbj+qaBMnpiYTsyCnyNV+ru3dmVgVOKPoQ0BdWj9CVZ/oa+2c
Ny/Cz0t6ylw1nyOZvdmXp/rLVBIhoP0BDIeeR45fvjqcPGS2UVPxHT5Jmh5q9P345GbWGyqTjVZY
lR4qGPKeME2RZ02VSHVetcaDxaSExwjaBevjEQX7LZXoCLWBvR5W6Tjdu3h7C5qwDIt49bTdiPvM
SOtTR7qlxjj+uH5s/rEu7i0dQIdcGqP3sUZSCEQfGpabCpJkAYdKm/GZuCpNG/TNbQBpLUSPce0y
E6jxG8hWX87gMnNaQn/8T6F70O/5ChjtfO2CCLWFl3t/wiY9AozTVS6L/ETLNdCakngPuXNab4LN
WmcYdyOwWZqxScMv0s7LGrGkOJw8ro7BNp1xqbCCm/r1DTgIK45NkHNmZAR/bQIInjcce/N1VsIi
brOTo6oV5bLgci+pUlcFCQ5RL5NMIBo/M7mZcAOHOq5itSPBovW7kihnaCpAq/j2OF6ITEeOF+/R
wsYTh2fWN3TlQ+oDkwdO7sbg8J7Nv2oS+iXxc5hiQ5S9pnnlg3QS7FR5UMI3WQy2faIT0Y0lhead
qT5qxC0AsUK3K1jsr8LVznz+/2uL0MLvBXCNzO4/cTTboCqNsEoMWBE/jZ1SdahdhFlwZb3cWWbf
wuPpOke9wZtqynsVGUjJF2c8TuhNoscj3YhrXryY/AYbIt7vcg5HXczuh/G/crlXk0K6QCwH1TRh
DWo0zA2oEuSN06mIljEe2sCBzfxi6NMLAYMx4WIWxhV7jbP4hXhucB97U0TPs+90bTmOTUc1lZ7w
2zpkXHprXQ4U+0hBdq1EefTTb+ss95pnM9Tm566TjnY2Jg1CCwze4AETXtgwMte5r89RzuEx3eUj
1zQ641bJOF+VAtamO22PjtZkGE69QGdAHdmVCQ61UwXSQAqgLrILGY84KpB7GMWlLwzpyao6elq0
hc1pLig8R3Ype50GMQP6IKjz/2Ck6x668r/uQf39iX75GTl4Q+5BxLUxmHbtXJw3NEx4bBw/8hww
I6bWFqpriWvlDPuM/EEJnbrqET2Ur6UKgdPml48M62Me0iIbPrGy7gMhFwDlNupKFzNHqkORMoql
FAubm7V20pHlJwBo6sxGQTfxtyDeInPr686N7HdcTuX3iOjZe2a6+9/griICNGMd+QDqii0wDZFO
b50kBeW1naV2cUCbGyhK/HoEc+HHhDqeJdKBHsSzy8/G+VUeV7YQUTI6eCZ4DPGHJkGpbPXomcbo
ppiWotljIb2j8aERFyJ3+OsnG673A6QqqQ2OBYmHYMv2IBH+VMINSkkKDIbznjnexc8tn8eBaiha
gTYlRrjYs+nxlHTI6r9JI+8TAtqEmhUQI8RO/haGYFKisysnZrZFY9dgukp+WasIHjiW4YTlfSZS
+ER0+SlbhHYJNY2DfQC8ZVZPbFZJdUAwjXevfaR4UphmYkTJMwre6E0wogyLkJHssfowfw+O8fYS
SwzCCF0Y0yKlWysmIas1J9p+gFyPzD05Z4mI29ykoPbGEyKxaQsEKzJUYpivERnlb0OxgU0geLzg
v8mfw8ovXsfCcxjApPQZPEcCe2vJPPE0ihp0+Q9c2SkNNqH3TH4M0Pz8B7JTHcG7R2YIYLj+dE1u
eZF1D8ksavbA8fX4G5IAQ7YhZ0dTUrboeLxzFu66XOHvK8G20nNA15U1xcGy10B29X4LWcE9hFgd
YsZrR00m6Vq1DFXq70im5RP3NNMz8LlGm0Z3YEZoS5JfK7LQRRtRh1b9vrYKZCEPbbW+heWz2GeI
ZDuHermfj51K3YQ9LrnF1K2UGtE6oOGGEGMcnxhaTaLi4N4NvMJXuMfaoJ8qzgmyvyojTV9Wbki8
YCIzXipbb7nPLnmtInGZb70xlAGqFdLO/+wg1Ip4FAXztXLs01itI+8B4LZfIeKhCISQox7aPtVI
ifXG2b37JnIJ2WSLNNMHvW+0gC/L9mqjaEWTLftQTkmy/nGW0T/BS+WlXpfZfsekUwmtbJW8mIX4
Rh7nKycbMLcCH1INChlqwCEebSiMf5ZNsoej+k3OGWkxNwwigSPeN56qqGZ/LsUL/uaFiCMVuK78
RsK6tAv0J/zjMykzQawB874PWLWSpJsP8jJfHCtTvVKx94IKOGOXlZnz2lbD6s+0uYu2VYggkQ/x
Y6P8JYF+e1Cg/vy2gaZVi39EHsFItoMvg5dXGA8+K+0C5zPbuJvTYUxlzE+inXbumRSTmKV+NYI7
kMoSexBGcsPzsoJsyQ3uv+9kQjwyClxk/gLVhu9fqrb2EJcokhXqq9a9Z3JWumtJlZhqjHZu4QKo
5gFe4SSIFBmWZY/H6Bdz8zReotG/xSMrFQwU0+w8rIz2lJvOuB0/9Ay6YfPEZ+agiLSdcKFiGU2g
Kf5D8s9d2JbTLFSeazwChoIWZP2Xqqo5d1z4MhN6+txHCvg8jSUd5NC1x5PSaM3TiNLfHT1YlaT3
VtKUI3oOwezxk1ksu/ngOfarS44c1hSV2cQgJ3kJn9buuo5vgI9aQei5tel/oYkYiHHFXxloEsrM
jFd0RUGBM3IbZlJl5qNl2T1u7fs/N2LjKdCSpSAxNCXoVrs4K8obzzF6p8RUYeeHzMsGwTGI7Ehu
XUUzJ4cU3DG11dBBiIe63ZHf3dfBC7qXFBgcdICzV8UrsborPK9Jo0+7SsPii29tSrLL2n28KOG9
nDPP1wL6fcYNM/0cP+1rAScoq4tZ1qaOYqhVE8AbdeJdVfqhniCwnOVhqSR6JAwKuuYy0U4NlNrJ
FMFIEGuLoLoEu501vK1a9xFpO7S9jaVAbzRgxoOc36jcyI38AWNzfQk/O+xQzM12L1lNXPt+pdBQ
WkbqumE+lctudcxWm6y+u3qCLF2IcT+gJET54K+rvxji1K8tbSPzTQduoZH6m8BPLu2pS3hCYkeW
JUx4N8ukuuOOnx9TN6eRfFs+yyclnsc6YG7Gts0hkJL7hb99AFVXZVgqClvnWROT7ODfZzQwxyM4
EzUdOoBxJW4scFHBQ5yge/2dhbj6+uLtjDTaZt+beiJt1iSIRNZibsSySWvf4PPWo/EnG3gs1VCw
JJpBP+zSJoX8Fx2lk2hoshamYPvZ9+/FKGm2XK19v4cth48f+AOGRBEgqUQf30B6Fx4flZwDTEOs
Banr5eEYpdeuH2waQpMDxHa5xoQ3fFQKIprubUf4J7rGg+mu0qBDYWxT5ZsB9tlEZD68DKCTQcz+
P+X4FBRS0540DvE4O5q9IcM1AavN7BtheQVhbl1Vv68+1pPbs+W7XE4uVpBCoxFCnr6h9Vts6ob9
QLwyPxUR9qmfBEm/yDY0adTaCe5Nj7q266FXlZpqWlbpXElTTrShVmRIHjep87FIWXyBAiDGQhZC
PeaITlO6uYZSktVMOd+2kujp5JY7AIQQ7QNjpqU47T/1mToNGWULBMx/0tN6PJnavg40psd9wD7X
Yv4+RymxUiG0uKezqdg7u4RCJie5PjDLwbPb4QgB+PZL5f1dPhD/JoAtUkabmM/o0ww1suxK/lx0
Ui3WUX7rrE+N+4Nr8O45B00MIB8EBoMNJPuUXeWrW7TheBtLXB/wvIjyDjq1S8JD8jKrfsLYW3bk
kTUqGOkdQCrUhQ3zgJj8n6muukGIQptVvLO5oibBf8Oik578CXQ+UXW0yMjKniF/qSzrICMrUf5G
UbsB2X1unlzPICUezkLIdzX4PFfQK3uuS7e2i1PNeESSw3JBbb9YrHLVGQJjZ/S7WgUpTrQUEjyz
DYCdEUNSE+K3VsVOduBdGv9xjm/8IGocb/L8IPy3EceWX5MAgSXWbPPZragTkuzEgyvsC9Zn1RV3
hRJlRAh6llRv2hbTY9P8Oyfl+N906rmvPVrvtwh4AbAVmPAOY++rIuZPKFqFqMWNGejbMQBmaxie
vWo/ZiiDiy6SkpvtETACsYvOmabVebmVM974qOESGwnq5PgyfRt3F1NhIjGj2jrVZ2ECypB3igQw
sTquMFH4Sm41FshFYMSUBpj+NoNPhXuzN8xKKxWUK1SGYFQOMkRXtukPDG4C8II0Kvk9RiWQGjHb
MbMe6g8kjenjMMwF57/KwXOgXhUk9tNzNT8ZkbXRHXVU1SU3XiKOhh6nuwYaWZ10x6SOC5V0o0VJ
dr4zkgFJnHbN1Iyeois7hJ5P85ABY+nBzPMQQQ9G7wxyBHMFi5nbq5zegHL/7A1NUGq6GxlP1qV+
5eBHnhuFWRLzzlvLDvXsUhwCF2ybBIijiVTb8vtH/Tuoc+koely4yTXHrfnKkNFG5kgpb5vRu/mG
F8wVjFEwvd72cQVU3vexcP7CLO1bW0J6aKwS+eTj3m4DKiUZAxzSjS2mQziMu8AwfsT4B8EFE0b8
NcSG71/SC8zo64F8e77vsQRolemoFz/M/NyVuCTX/xTBk5pWTppbiGSbE3cuQ5GrEtGxnYlT87Ds
F5rvyI5P/jhey3JEqCcqpQ+JOHurDII/jrMLjfg1cugVVfht+d+S8jp2071Zp0e5pAED7bgVmR8S
OE0LpLVIe/8t3FJnp+pE+6BcYqe3WBRq9ve0bLWL6mv1+jWTaLlWH4pFbz58toBjLTnOxu8vikjD
1QMs+ojnEfyNGG7/j0K0/b3voHRiZ7qgfGo5QaQBZDKQPSBIDsJTd17+UilQR3qZFgpRdbOPGpE1
mcynqNdzp/xw4dD0/YgIA96AL4iriKv/sCeVvWI+BJb5V0ENmsKrbyFThzsaD4jOHzkip+6HtwND
+vqZ2ZE2ONIHsQ4lhWMt59gH51Ch9BpQdvLBPyW/RkcrEoqlNIRXiW1RwWYC+PlITXAAtTgOkIUm
pDWc+gPxPxlqvLn09y/B3eJmQgh0Y9CCOubX8wwHmZMwTgbkh08QtIzZBFKLbcQ+2wi+Jq4QSSRf
LtrUJgH3HRe3NosgXujnO+3or/k/flWfQmp4dzhl30CGUwpIsQjcFsUABKmQ45J+MsBL9ZUuSqLL
7AM8RYAPMyB2tQpUa4qHxHjJGTjF9SKWyHZpxRkWKhUkLYcdY1StyTC58QIaWsk0JfU6EH0JL8bE
QpDJIyGuqCfuwXdupRhT53JrC6SDkOX5C4qfXhj8garbfyvRgAReO/pUorT2nZiVCe4A18fYmt+0
rR3PzwkvCMCOwbI+94doVq6IGn7Ul9lQszR7y3TaFk9woWB9WPekVlVApuu5mtmxl1ixq/PxJHo7
ma+uIUhL/w0Pll5rh/3QMRjAD68Sw/m2eNvBIJ0SBQ9k33E6Mnsf8AsshAkQ1I0DLONT6TmSwBzN
03xQx99aflNe/mJrccRWHMXMtNYqT9qzZeQGaHMIV7/WAMSg+QJsWN5B6xg7OHaaokcfiHkuqzNw
JQo1kA9kUv4jO78i8rtx5YC9q/sJQNlwY2T8/rsOeHHN7VZ/yCM+KcIa6rRFLb+EpIgMgo7Maavv
V2KcFvL9pZv6xNSfJHw1rANFqelPVees/56Lh/BFk8XZrQJVatbPRJmyqZM68VtN8l6h2uKOy9Qs
nRZmixXxxniSpjeFcl79DtK1pNXnE6CEzwsBipLnoZylPbeD4wt1QEUuEGJ+2bX6edmKOiWVLXPV
0FxdqKqVXu1+JVhlytfEd+pzmB/BKwVB+VvHWMlGj1Px8tMzTFYTKpYCeNiU6h/P3mTSv1mSA1SA
s0IQesOnV8TBa2zR/7l01KUnmMFUWgDKGJEDxI60thEtuVbewSTno5iGV3cNIE9uTDnS5I2//90N
N6mCdTthyiPn1yQW6bJisilT9Sc3RBC6tzi99NRyr2m6/TuFxO35pjbPta0MpMPpVU3lzIHbJlDZ
1EuFzTabb9atRK8C29tmZpYS6RbWboRaadZrDu0ixZpjAFzfNMAyCdVL0nIZDEAVNFb4yEfLwIab
O75LMCJhH1gs+iNpiFbEdXcUM4TgLNyQjZB/NCjtzAzW480tPpEbhsMmzpHYojLdBK2pJWfqxwIY
hnDyaxqUgMCxIN3w0l430m1N1D96rLKJkg6lIxjadEfmHPyKU5KQZSQqoDIA21wuX6rvL4kd+0UM
gsgz0e0ZiwalE+lhbqD/pqpCnsS2X8gpDBodTNTab2t+e9ZjceA102PU0/krOxJfJRK2xfl0NKo+
Zdkwy0PESrAfCf3KgLW9o3iU/pZcyewpYecOpet2oUyHMLLrlrOpfIszgPvJ+CSXQDmhCSK/jmmo
q3wClwxx+fKTkGz8vbu0Lilo0h75O9ElpASz9A8Gnlsc4fgKGI4dNz7zfbDmSE8f7pnNnEHWBxIV
X8lbZPefQOyVcl2Lj5Xh5Oa2JFI0T889+2iS8CTtoZCey/2cQiSE8+NuGHILgh7+hA+cozd16fqm
FkaDL43ClBqKIDeho5WLuBiWp7AbYx4QfuyZh11HBPw8AyVKYzBjp4tfpgQqIvWE7C1IoeA9uhH0
Cdg/JSwgI8vUSB+hMuGdcSPLWtkrF+Qb4DXSGKPDBiv0FulqcEwuNcCJsE4xMAEXTmcZZKSZrOZt
BklTFeKXZsBw3dPzNt99ryQPYT+dETBSrcj/WrDc//dNtjcfyNX4bISP24H7IwTsTXAAdH4bdatt
g5uK3Tq4Jh0a6XuZ0uO6z7WYvPNGfvGwjNEVn3IucNp/plGNSu8q9Yxap3l0ja0TVWxr1/9MV9Vq
9+rrNAoUMfExW4x11TLfKO4je9MpE4XgUo1eY0Vvh0c4CHGB6MEe1/+/LBAV7wXc80bhrsZt3EL/
7kxApnRN7BE192l/Uu/nJXaAn1QI3XC082xdto0mpwyWcPlpt9hi0zNhExJMfSuKq1DeCloP+huJ
w2AaI2VyDOOA4wApmJJL0jcRq3EHfiV6rTZ2ua7Jiy8Aofx1x4EVpX0AC8QDkpIgah35t9Uq0+lm
cGMD9X6PdyBBnmsmnLuuPsOiIYD/xbRZOxaJ+QvG+goh2hn2w5rQL08SoNgFN0p6PKUdpusR66bs
Y8rSPjgKocEf29MaCPccghQheDvNND1LOXYXXf9AZRk/ogKIb3hLOYzCE8EE+B+UhaxxkXfW0xDc
ZPX57QbL3sIJ0cgRPtbEwCdSVPj6LkIynxq5FqBrkS0WoD+3HJEAIwin5vMFlkVWHU9bf6T5TQ0Z
ZggBBCwt0cM/46TGOSW5eoxQXMSUOkWJkziUVWRME/4cHYKCNWcBjldWscbJT+pJ0KN9ND9LDX74
/BJMmtD6m4WIv6QEsiklMwQpHgMMTyvR7ftdU3X5shxzQPeOMB/SDEiG7/qEag410vF+uxQM+ooJ
Qh2XWGlbI4NL0xZ7moC8SXN/6SWsCTie6io4mtJD1l8M4Pffc63nZ7tbqjE/PrYL7DgZKgKQJzRE
jR2+klsymcpKPL6eApuk029+6Bseaj42q3Dd3IGvTQvGQ0bQ12aqi+C/K45G4xHDtBs6QjKEn19n
4ohbt2Lo3oa5FqlFFUqfsGL0TU+pHZ1TBAMzvJuiOU8qx/u6eb5mE1uUzbw10Y5tx6PV5NL+nZeI
TcaZu64OO+BBHk6jfWuvwAkMxE1PLhwb/Hb1EWaCZfntxs+B2MBGGJgyRt+l17+8MvuQlFF5mmL9
ljvv4htSf7otptnzndZ38OpEDMw6IBSmvP1yIPyO4ACFMa/Ra2cf31833dzPvRkh+oTrNU70RuMj
DzzxpCAPIdvFjbQylSUNNFuDPhwFT6gLgPOQpWmbwegWUKcrRVW3Tvi2/7eIrRe6CS6v58lNqQRL
RWWsefnsbzhunFxzIM2nYYiMiYaqcw/FtX0JlvNiKnFQW+MaJfyBTSibmDEH8NJmoDE6+UayBt6U
qs6pZCGP0PjTXrUCRkrJldm0MDLcL6H+MClJkOZfYWQB8ZQp166zDbfqL6Q3IOBsbZMiz1jL6rFZ
Gg4R/H5cMKADgAJ+g0wtg2En9beuSv1uZdWFePtPTrgwo2vVr6/wgNXOnDtmhbNT3U0vwn4MFrOq
qSxwHjpSfVwOh7Th/vAmuBu9P/wN11P6bzy4gnARoduaZD1W9tEL3WaxpqwBxiQ0LgGxndl7io71
O5pnh9wntpcE8LrlcqU9iTKzX2DIJgbHtXmU/2ZJJaAMB5/QHErYqD6vMXg0f8q+4E/RuA2PRbQb
ZMER+QBsP8YD3R3yqZIseT/nc129LOYwtXY6k4IyUSglNe51XqDlaHM0FNWkLokF/nJQxyjwQyqA
WC5bUpYSlKtGHE/IejA4Qk2A5xaGHZKVIr3wRbGxtQdkv9XpKuEscDzkSIBJJA3Blugie8wXNgkt
r9Gq7tEhdSaszG4HqgMerTioSp3xPGhIQtSz2h2RQHOmTXHbrmBvLMP8GX0mitNOscPIUO4IwnBO
UdvcnpcydWU2kLCnCSYUyLidQKsnsFSItDFkGuvAKp7a39SVnV2K0ZnBhL7XPX6a9fJcSWXKTjqh
fCpcCizfAYtKfrErPSFyhIvoVasVH3gy+XDCANfTWYYyPnMVPcDUv8UWk1/ljFUMMhogOftof8gA
agZ0UcQaLpDLUifHESjWFA5+EGcc2xi2h5VCgmlJJOkYpqY/UoxdaRIIT9hJDv6rYiJa8oewVzJE
ErBQoB/56b38Z2Ie+DjwzRnMC2KES75B2u9xENZqxJ9qLLv+FPbaIAK4PMVV+LpQscpkyv8ehYzc
SDUpCvN6tPv7D/LFX90Kp4gweHHON7Wso0DAa1s5uDhXiCNcxnoHhQb1BqpOfE+sFfZYwmR3g4yi
2GjKTLKyIG1kzCV2rAVJF0Pmuiuu61lNqDQlqBDRTarrAN7ZeIi1GV75GUgA1Q145FI3hq2ppAHg
mF3gs83TyEBwKiSRftUoXZgc3GxE3AaZehXHqKC0JqkJ55vYdjf7BkoRL7Mvr1iiNuVvX5MN36yG
BulRITTaxipDNATMg45vjuDFqSk2CzE9SmlJ1DrHKVMV4q/sVb3A/vstpzI2I6zlczQj5d4oD1o9
QkppiaZn3kOicZ8VhX4XiDJ9SRZpYC6joRP++9Evm+KUPqbJKEVK9qk+f9icodWrXch5XrA/6TUx
1gWLhbvovLXphlDq1OTZkffgb71b6NYBLVxr+LMiI+KC9juM3VT1TrA6cIbl0RtzsAEpimtAx6V7
dIBxz5jW8R3+MX0omObveH6lWH6yxSQR6SdbIb+ondroFZycuy86Rub56auW0vfB0nqOSjlh4r2D
1TpCnBlVkYpGPjYDS5Rgc39SKZXRNdh6AtS/dWLm1lebwynfHO1T7SV4eIFaKKFn7ShQpDAVcL3U
lSM5m0D33jQKKesEFMOcImNy+Nw3+D1Xk1pImFbaidx354jDhpysGRKl2FwLNnHln9VbfZp4A6Dv
LsuR34/bIJuBLFZ+JMj7rZKcxwt3Q/5YDaAOW3Vd8vEMH7Z6dUiRkuJEihz+xBGzKmBX9/xLUHoQ
ylkOH17cXtaiJmn1RHE8vOCqVKCilm+HUSUi+NyI5mSqHvjg3K0HjZj5Z30QHHtptJGVKTqMuxKU
7JUHHebywczSgu7b7k5FxXiHBoTR6Y0w/TqygstTUjzC/U+b2snyJYv13DAkfdVngacjX2NM8MrK
diY/HRUZxv7awvBBJnKMUgUR8ZP/+oYI9D5wDYWnLeO3/zW9JaDff/LJoi9UeV+j/1Ysgqdl/N40
mhN4O/wmaLWEvCRwmX3q0/ftZGJmSQJDCwK9T6YHrIZwtW5mRT33tShUYL/mkUZ1tHX/nqcly1iz
8WyG3v3mXBtyGn0xR+/zFKmGdNr5qddbBdQVMRgIAF1H+AjDu/X7Qp/R4H2c5VR7cwbq4XbOS8qB
kqYZYyWSqqsJKeLel4/lfFs9WG3dTCiGiwNYTIP48ETbSfQQZ9UEjpdQLCZv70snCikIwdOoDjTe
+stVGkylum52yV9HhHkI7JkqXj2284z34cCfsHmSLgBwSr289XolkQpTFXSOJevwZnrjPh9oSX8c
BdZ++0UCQKEGLXY4XXmKy6q/Hv430F25oI0BpkdqYVdNsg/IH5PAjAkvdO1hTCL8iG3/RlqO004D
+KXbYPFDzgy1lPIWpb6yf4OsidTKP5rp8aSgctIQWkHIm09DwXasfxKM3ma5afYasaRl8qNAUBmw
AVX5tpe/eyHqIyRmy5KRUPohbi1r9HFKuacD0mLjOzQFF3BuEZwgnfeojteNkveSMzqdrcSfE+Yk
3OkZ5eYrbBh3vlppyfNfEzscMZhCAYdBgQWbQkitmAIkWfuC6xeurr3oqDQ8WtByh0xjvQyxiYXe
4f4j4itjeh91rd+zj4cQ2xe5eDj0wckVj/lsWha26J124DLoZBhLIgxZRVAQt2JjQhd9bA9KAbkt
v02Vt/v5ws8VgB+uYIJK5FDwm6gae/3T/enuXaITK/VfoioXcSPqfd3/S/9LqNClf2j4YQ7y+fWy
GEtLhtkFjU2EQoWuevhBpiKWM352HoxvvO5k/caXYeqsZGJjTQGsonKmoPyCTr9pnJ51bv9kcVWp
DqLe/J5agbHocGt5V+ghavgRXxYQqbZ8daDW2kSau8/utwbV7WAq3jo2mWsODPzZTCh/krrooFp8
ZOnmELr56JT/UyvXpY35jH5/56wt83mbJwUySuk0Xx4EFUDxUIG4DeOdLlsrw78poj/E6BGEWprP
BQLW9O/sasEGxE6eqaOBWFdDHsTtLIGUcu9EEHgQpg6tLT/OWVbDH9bE3bEHMmEyJmw3LuK/bdib
YR5OeeA2oyf18WIh9i2D2s/gf6cCxQ2y4srFyOVPZj2Mqq0CZC7LqrPKDJSo6NR1kkBGOqPwjuix
kfjK1KPjRIIfycdFiv9/r5pfxq8vFRGOME171lIc2EYE+UA7HM9ZM7xMbZJKm551pyfGBFDB4bKd
b6xbT7EI9PavA9iT0yLEkf7pjH6H+hFOEnMeiIoReCF9s4hMZpGmZPMPNa/hkbwXt8UNEzYUMYPZ
V/fx4g3c3HNb0kmh1mT0sSkA46FbYCZhsVJl6EWnMzeaYl0wLw4G50ID+vz25stUE/7Lmhw+qFsx
4BH35ScU2pnjjW7phVD3StAQ2UxD1S+3CtdztkpQVYh9tSWWlAb/d7DrnL2MbJuaZiPXVu//87ol
RNJ3kvvGHw6cRoJvQ4/0zMfztaKQbr6glBKXdZsKeUAqeZTQBJ98kZiZ+ZAAG+MypzjoSKk0COOU
8/VrmRS5Bp/8GHqeNorNswHMkUkC28fqH34OL2XaJNGeOOUlQJWOaZpJmnCwQMyk1tbbv6jaCNLr
svxJ5pd2vCv8Mg78p2KjHCh1pUHJGjN5uDFGSOsL7Xua04pnlTfUrbw4NcO1NfwRFqCBFsBcAZSL
Ah5zwleDqdfncomjIaUddPkXfOyyRNHi5A+8Z3B8d6y9I4IlCXEU3kiNXxzoesfuzIkDj1U2krUS
4rFt0V+LJeavYti4lCJP1/VffJWK/Dby50ko1WVkQblQegwf27/BrWeWePm1m4ux+4bd8pagBlm2
LaFN8U5b2Gyn4EF+asPeYRtsJ7SDVhXoXAIUIULfvB2YEAj9yMkEvM2ZSbz/yBqrebrXLW4KQ3j2
x0wA2Yb1NCwV/8sfizThUvYucQNJXpJoRPv7qEM4KVy3ZQKmmBgS5QfEFu46rK5ekZ1lmJtH6Tgm
MjMR2UpqToUVvL8tqcn2OK/NP5v372ru0kojI+xDqCZqoVWQTPITHLkuCL9WZTcjgQcreiVmCNQj
FxnifMFkDh46Dc5vQMpB9yZ8ndLnXmItmjdXESZmmyI4f5MtJG1wBfrEpUE9e71BgluBqZ5xNdsr
IUfBbTfZsJHaTN0a/uMV/1s/Mhv98OsEX3lJBKUzOjhGVoE8xfjkxH8yU2odjAOtCx7KMSI2wpka
UcSx3eQ5FLGdryKFLh5RUQRiIjqZG9bItzoTYB9/OE/8RcvjHBII2YJcT98PF8zCh24nhhQYdrRb
ybt9am8CXKm+5OSb4u6l8plmyHxkfzjHxTw3lR9l7vu0uNhKlM8+I2GNlatYm/WcGrUBPQQP/ge5
4Fkc/wajlBKPKvnKAf25Y9dC8btXMSvJPdGW47P78mxUHTdxM2bbSIEkJogZTAYdUMGap4RoYYMU
E6RbVmbBXbTuh4RKfV31vIE79rqtpt6Itfrkg4gmCFrIBVoFIUOOdAViEW7IqQU6TJUJsqbXHCS0
9Tx0gBYss+cZmfkOCybl2teQApLqSoqnH72vAgZCoU7LLi20is5mcZ7VuyIcUc4VPxWF6cG1ZwGU
ssFnaohk8/E1lQ9xO2zTsg91ATIv8JhcyzJrTGGa5fNjDdGFCDX4OqvScCYRAb+KwBzp9OWcQlMA
Hw3yFhYGLzwzIZJQWYFBIq2i3JrbtHLiTFFLsnsXfdxbrgCizqjW66aeE4ijoK0DX+2Y4sJLw985
7IjoAczpKmn/FD6bvRE5eB6sF9rjT/WT4As7ZHEvKcU1zGBhH6yECfzky+jq6HMGOGMQfg5DzVXv
RkLmzgAlXsdRdqpjLu9LWU0FfMFEEW1PR6UG2hxPk1olBwm6m/JBgVsQB78OJk44N0BZ1fGXz7Z3
z60A3wtcroGe31/YWZ3SaC9lBhDhGTPHOTGVLXPDvGi8/IesRTZfklSf7PLteyHy1wziDFXMZ/E3
yB+bqM7e5XgAicNVu7g2gLeHGB7MBDEt4zWYLT0SGbrhsfawkilr4MXJKcyjQ6gGBbfFeDNotghp
0HBfVMRgLuz2vTXAronVwCRTAPqg2k5HjSEs6r5tHTs37T+1owwnIerp4ctERIw3sMry/XseQ9NV
x3bzWCjGzlFGEpoB/JtxFRH6ppHUKwpzwEKVJb2hW5NNkINNr8bkkD9jInARq83sLIQsJ82ifPp7
oYHlUjPlcak5mAVZKC+/xCo/vqcDFwwuYQNQS8Te5OCGSlvGPx5d7kVWSdWllY19lrASYppYEcM2
PXhoIvNtPAtmO61jyfUXwk/YDkv+eK8ycCbv7an83L8z084JLh5RKiBESYj2HExtxr22wJv+L+Mp
gP2ohGsQ3Rud6dHCjT+MdedWVAGfKjtwb3vRBrPKyYxT0ngUBEGggLfRSI7YJcC8u+DsjcXn8pqw
sK6SL6hUD8tTNBJlnH88zpCT4dRGqSItOUeSYnzp6MqWPCDs7b5ALoUs5MTjXtYZIMhaleVyG5pH
2cevKFVnc1bR7HMSy3T8xX/cyj3tbAKI5dVwq7Imj12ge1GxckJ6z420xUYzH3n5XpJw013Ai7yL
p5to7WrbqQSPNLdAcuPCseglnd6hZwn9jojYkS8mu2rQIjUqXhUZ/DBRUBk9RijDH0miLSA3rJ87
p9m7VAELpbgfv3BNFPqKXulZJNJ3bWGE55pESeLkU8PqmthPRHffWk4jT04tCLcaq1hPKVVrx2Hr
MAG0tH4jRDRKo4q13ahm2uOB4TEp88SACJKZnuxg3xpxryz4dBR1w+QvTwtjvMAZDxQGmcK2+9g0
H4Z6TsIuR9/g7ZiA0172Iiwt6ZACjbzK6eIK1C44VyQexjKXBKteEmW3AYUzfaS7aQKxcr1u6/EY
HtwfXdV3coogHzyObYRlcQIW71v86WFfrzbgZnzqZsCOHHlIWhpHhktr9i0IuVkmcLoQY+BdHMWJ
w1oX2A2wtAzD4t7R9/bTlKv+2YmGCuoUYEiYCNCo3TafMaR7mjmurf8n+n02QEKqyvhyBnH201nW
dt5/bFIZ1/i5ki65VZdtuorQQOIirsmFbbtJ+dQX9n/lXg8gX27ItnB/3sdzlRg0OUCuia6R/tsq
pBi3HjKSZ4r3wg9FtbQ8skVY/7nbhLOHi5j3E1CENQwO0Wxv1V0k5koCFieNsPmmrbOsK3Ujm+7C
PD8ElLhYDstXHN0mhLcna9FaN27FcdKB43gYUC2WVJqMY/aWmmUkASMvWcmAMdVKmtYItVxSj4CC
7U7lQjzpJ4iVBfnRe9WLcSPtgVJDyYs7pj0cpb7LM9/sbIEGTLU+37HrRjCWaNahg8g7Kv9A1/Ca
i6M3Fd1+G2JXFEKBPpMH1w/O566diKiMqJhDUIui4R6wFkCFqB4dE1Eghea82nKJA6J49efVIWnP
VCYnlFjdQ9XtMmYH9GrhVxXcv3AVn3f7rxnOhRxeTER51DG6U4821IgV0XFAoW10ANxUOx6l/V3M
CFrFk92/Q19Fx3L69Qu0/457JV+yvA90EqPWEjzfu7i0ZMtmsliLNVIkOgq86SsjdFyhy0I+n8ci
5177s9HhiknV8plBpw6ta+S5ZsHrs2jFKcWI97HC9zWM4bkoMrmOeXpBjYM5w7mdql+vUZ3l75Fg
EeFFX4I7XqFmerJRuox1I2K9gecqv3HGJ37EVt/3qW/UzAVSdwjOD9X60/m71lLDe5CHzE8pXXht
t3gx+46mdanVEwDYX+hK+To8IjH7MmZkqMTBKiBjz/gnR4vliHE6YTIDKbcJ8YNT/DXywFIhJY14
Ec5QLAbdg07X+PPwRILA1E7KY+AfRaTFdumEIh27BXbTFfqO7iaDQqxkr10SfDaOZnF7E0fHC8hE
jy0qg374GLizicMdLCEkSA6TZoGHYkJYsyywb1V3DuVMKXvHmiUNXaLk1E4EfO2JcGpqziDUavJJ
bzEk8zs8XhJ53EpXfk7hGW/CBYodaY/Ju39U9lwEzs9HX6nObbDWYnO92yp1HcfBxURkNra9Y8C4
JnGzeaQRGGoHvo/zpR2slAdlRNyc5uBZ9K9Ep6Pe3ncQpYFUylq4dMPXknBsYl2U4cPROM1oy+Ax
YEmUvQ4LCBcldCbjgGX+dvC1/Hk+FE6nl8UlSE2mzN5BDFgCmTQj7NZkpxiex8Mh3wfcgnE1ZRXn
yKNREs0A57CPFqmtePM4cTXG8rDochu7D0LJtRPMlShf10yZ3v+Dz//0c/FDACDVU0vezEDJRVS3
xoFTEer+I8TLRUu+BpdMt1CGTvDHhC7InxnarrP5iB0eFlU0xyPnRETbHnm+ljst2qNvSuQjJdIq
adSoT6J5YxM3NSxqCTYv5PUGwhKsLu4mV74hxKuLk9njGFj+ZwF0hHxQrAZCafF88N2YtakSyb33
XnfjwnFRXoN6GdXaltEJwRQFrLRQbl3IV1c5SBAs5FvvhPMwSXAjrVuYY93wGcWZgDiMHi1zROtS
KDfnfCJ8ElmbfkIMumQJNJoOBUa2a5bPTxg/CZhE2a/u8xKqrWwSEWttbWEZ+cVKINmSsg55yEfH
lYpH6O4HCa9piNuw6ZFFdEj4QiomEk0TAHbMoWtbUs1kW/WGysHY+wXC9Lv+mSaysi6pV0a5Wr5B
X4p61BN61Hm51JEKRGEtUQ995wZnHbDoikkTgBNHHXTsgP9uD3m+FNXOBWc8/77ZgsSZL3hmAY6G
sGnkV31aC3U8R/YERPbRwAj4LCfDiQ3eUmD2bT0Cti/Px1W9nbW2B/jWNt3VoBJ2DGR6A+csOcER
WOAqJ2BK/nyyJJ2+JMlgtIqgGcgjy3ZzKoC5FN/1fuTS22RQXbNQKNrgDq8w0em0uJ8/GddSx3N4
subYU8gDbrB+8TQxxZO/LN814Mqi7NmpogKYnTogZpdE5hiuxc1F/i06suLaL9UjubiIVuLWTTK0
xXFzmv9iFSEyAWyB0WtgW77mCoKsR2tD8KhfAk2jH6frPlBIC4N1LqaAZhu+82DlW9fv0/t30k8i
+ziL/4fhwm5Tsj23QB2bjyal2KhAiTs3s5To0j7kOtA/5ppy431K440zPjADDCD3m+gzme/2q34A
8K/vQ0sBFyxWGc57RcdsXeRcXaezBX0J3o4BgWFikBBLH7W+eVZC+1qrO81ZHxm+CFqwCaG/oXed
deTG/67DNH4J1Q8bjk8n+0IWUV3myCwOaJtByNbm4aJX5OSrEpXu9+udqNNlOWBbolxgWPZ4L1DO
GlGt88CC0MBMAqFfn4WSkdxxSKT4xHMH3Ahy469fwh9ZviiaOYlpnojenTkZnQz/v66qUnJdS+G5
MzzAbXJUs7gqo1QiKE+wsHqbqsE4TstWUczxgou2GL25fflANeih2LDEFnoG0Qk2GPTMvxj9Zptp
tVEKG8SGmgDZXQJFab9o9AXql0n7qS35FluFT/h/tasMx9buJapUavjw9DfyN60Q7HQR/x0Al8Di
ipjtE1N0oFbw32HS+eJ7xvvB41xAsp3krDGfnH9DcmMRsSpaTyjVm2+8dSl2K8tWVmcLDq6My5bj
34ndwLmF/VrggEBw7eiIiO2BxCqSYK+sAZu5KaQu0SfxHfTqyC0lNZqcwSFsKBSeA6rbgsh1ePlN
AJIeIA7Q3C2ESFoAK3W1IbqpBGd8e10Lbi7ndJqIElK2/8U9cytTdIk6lugKIQlF0hnw8JtzvNAT
vDJqLV8P4rEZqKy5nGm4bZO+EoLBIaRAgYvGebh/TJqb35NWgbrvnTGFBWb4HHOh1U7+wwLRL42h
SULMLtTSYKCVYuXM4aaHt/ZXj8J8OZklrUozjtO8zLpn/3pG0f5mygfgIIz72cSTL2VjOTeZYarC
59F1bsCbbXiRGzQQTKhzp1nqHiZSHefDq+c+0josVMRYovkLSHlrvHE67exEPZS1mBGM+6hnawkZ
hO2MYVBEvKQ2sC+IwLRVgDBTK57MgKBqiA8deyMt3QdLDyqMD1kY3Jlrj2F3uWMrq9BxmQqhUiUp
sPXzTJDaqgumaRo0VzzGvNdR/lN2sr2lajShJ9GW+zWGyn6X7Nter9h0Hkntjqe2kQ/xCmApu72C
CJlel9GY29oGPbpfrTaC3+Ct1mHteH7OGfleP7fOO+g+AyWfo56UapsK2GVqq6/hfyOozQRIkjIb
qh+x/xzZFFIa59YYwPN737ThCYTwNUcTQpHaDUbR/ODUifE2Hwnj8mdiEhhzt07JxZUeO4vhZrTh
GH06jAVrP2YzN74EjRsDugO9ijiLDSlXmYx/1b7Wn1O2E/HgztfgzExGpiVFZ/Fio9lp1EvfDiYM
bhnUSIhYKmSgWPT8U0rHdXjnpO10JX54C4Sw0Ybizi9rCNIv0avb3uaekMgbKS0TozrSMjszBh0R
8NxSWjznEyAb8u9JoSTuWicAL/gfGcmMr5qhNr9ehFAdQDhPMWWP8013B9LLryG30CxZNZSRxWZW
pRamU2cWx2IOLx7xfeybWDElAXsuIVnMNUwCIPXr8NuKdiEyOOr82hHa69GJPDTKPfpm0g7fIXvY
+4f+p6THBf2f2MesjDIyKYKIj4bKsMo2w6iF3GWlmxEJK7BvM3n4ayASSq6KvSmzEXVpGnUgUYn1
jswWgZzQG5flKgZw5myt+n7XHEDS7s8rfeML0MXDVRSQGsNjtLiKZrrcBp08A4TuLo1Eizrkx1us
tYMBHQfdSsZQe/rM31aDyXMBYOy1rgUuIPkzSfBQYC9B2dWNBbuOoHlVN/sKfHZlwTgbVA==
`protect end_protected

